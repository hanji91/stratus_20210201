/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:13 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3784,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3850,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4000,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4017,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4033,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4059,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4784,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4850,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4866,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4921,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5000,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5017,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5059,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22921,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22987;
wire N10691,N10698,N10705,N10712,N10719,N10726,N10733 
	,N10740,N10747,N10754,N10761,N10768,N10775,N10782,N10789 
	,N10796,N10803,N10810,N10817,N10824,N10831,N10838,N10852 
	,N10901,N10941,N10946,N10951,N10956,N10961,N10966,N10971 
	,N10976,N10981,N10986,N10988,N10995,N11002,N11009,N11016 
	,N11023,N11030,N11037,N11044,N11051,N11058,N11065,N11072 
	,N11079,N11100,N11143,N11261,N11288,N11290,N11293,N11297 
	,N11299,N11304,N11360,N11368,N11372,N11377,N11399,N11401 
	,N11418,N11462,N11464,N11515,N11528,N11530,N11536,N11538 
	,N11547,N11554,N11556,N11563,N11565,N11572,N11574,N11580 
	,N11584,N11586,N11593,N11595,N11607,N11609,N11614,N11635 
	,N11646,N11658,N11665,N11684,N12025,N12031,N12063,N12074 
	,N12081,N12084,N12086,N12091,N12096,N12100,N12102,N12104 
	,N12110,N12112,N12119,N12123,N12147,N12417,N12418,N12419 
	,N12420,N12423,N12434,N12440,N12523,N12531,N12533,N12551 
	,N12555,N12573;
reg x_reg_23__retimed_I6694_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6694_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22628;
	end
assign N12147 = x_reg_23__retimed_I6694_QOUT;
reg x_reg_14__retimed_I6682_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6682_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7520;
	end
assign N12123 = x_reg_14__retimed_I6682_QOUT;
reg x_reg_10__retimed_I6680_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I6680_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7437;
	end
assign N12119 = x_reg_10__retimed_I6680_QOUT;
reg x_reg_23__retimed_I6677_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6677_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7738;
	end
assign N12112 = x_reg_23__retimed_I6677_QOUT;
reg x_reg_23__retimed_I6676_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6676_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7744;
	end
assign N12110 = x_reg_23__retimed_I6676_QOUT;
reg x_reg_22__retimed_I6674_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6674_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8329;
	end
assign N12104 = x_reg_22__retimed_I6674_QOUT;
reg x_reg_11__retimed_I6673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6673_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7530;
	end
assign N12102 = x_reg_11__retimed_I6673_QOUT;
reg x_reg_11__retimed_I6672_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6672_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450;
	end
assign N12100 = x_reg_11__retimed_I6672_QOUT;
reg x_reg_18__retimed_I6671_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I6671_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504;
	end
assign N12096 = x_reg_18__retimed_I6671_QOUT;
reg x_reg_20__retimed_I6669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6669_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7486;
	end
assign N12091 = x_reg_20__retimed_I6669_QOUT;
reg x_reg_22__retimed_I6667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6667_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7469;
	end
assign N12086 = x_reg_22__retimed_I6667_QOUT;
reg x_reg_22__retimed_I6666_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6666_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452;
	end
assign N12084 = x_reg_22__retimed_I6666_QOUT;
reg x_reg_19__retimed_I6665_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6665_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550;
	end
assign N12081 = x_reg_19__retimed_I6665_QOUT;
reg x_reg_23__retimed_I6662_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6662_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7506;
	end
assign N12074 = x_reg_23__retimed_I6662_QOUT;
reg x_reg_23__retimed_I6658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6658_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500;
	end
assign N12063 = x_reg_23__retimed_I6658_QOUT;
reg x_reg_11__retimed_I6642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6642_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7446;
	end
assign N12031 = x_reg_11__retimed_I6642_QOUT;
reg x_reg_23__retimed_I6639_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6639_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3];
	end
assign N12025 = x_reg_23__retimed_I6639_QOUT;
reg x_reg_23__retimed_I6493_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6493_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22622;
	end
assign N11684 = x_reg_23__retimed_I6493_QOUT;
reg x_reg_23__retimed_I6487_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6487_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22631;
	end
assign N11665 = x_reg_23__retimed_I6487_QOUT;
reg x_reg_23__retimed_I6484_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6484_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22637;
	end
assign N11658 = x_reg_23__retimed_I6484_QOUT;
reg x_reg_23__retimed_I6479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6479_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22612;
	end
assign N11646 = x_reg_23__retimed_I6479_QOUT;
reg x_reg_23__retimed_I6475_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6475_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47];
	end
assign N11635 = x_reg_23__retimed_I6475_QOUT;
reg x_reg_23__retimed_I6472_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6472_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854;
	end
assign N11614 = x_reg_23__retimed_I6472_QOUT;
reg x_reg_23__retimed_I6470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6470_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22871;
	end
assign N11609 = x_reg_23__retimed_I6470_QOUT;
reg x_reg_23__retimed_I6469_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6469_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22865;
	end
assign N11607 = x_reg_23__retimed_I6469_QOUT;
reg x_reg_23__retimed_I6464_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6464_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004;
	end
assign N11595 = x_reg_23__retimed_I6464_QOUT;
reg x_reg_23__retimed_I6463_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6463_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[6];
	end
assign N11593 = x_reg_23__retimed_I6463_QOUT;
reg x_reg_23__retimed_I6461_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6461_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991;
	end
assign N11586 = x_reg_23__retimed_I6461_QOUT;
reg x_reg_23__retimed_I6460_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6460_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[7];
	end
assign N11584 = x_reg_23__retimed_I6460_QOUT;
reg x_reg_23__retimed_I6459_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6459_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22677;
	end
assign N11580 = x_reg_23__retimed_I6459_QOUT;
reg x_reg_23__retimed_I6457_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6457_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[9];
	end
assign N11574 = x_reg_23__retimed_I6457_QOUT;
reg x_reg_23__retimed_I6456_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6456_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9];
	end
assign N11572 = x_reg_23__retimed_I6456_QOUT;
reg x_reg_23__retimed_I6454_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6454_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[1];
	end
assign N11565 = x_reg_23__retimed_I6454_QOUT;
reg x_reg_23__retimed_I6453_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6453_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1];
	end
assign N11563 = x_reg_23__retimed_I6453_QOUT;
reg x_reg_23__retimed_I6451_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6451_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[2];
	end
assign N11556 = x_reg_23__retimed_I6451_QOUT;
reg x_reg_23__retimed_I6450_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6450_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2];
	end
assign N11554 = x_reg_23__retimed_I6450_QOUT;
reg x_reg_23__retimed_I6448_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6448_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[3];
	end
assign N11547 = x_reg_23__retimed_I6448_QOUT;
reg x_reg_23__retimed_I6445_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6445_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22861;
	end
assign N11538 = x_reg_23__retimed_I6445_QOUT;
reg x_reg_23__retimed_I6444_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6444_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846;
	end
assign N11536 = x_reg_23__retimed_I6444_QOUT;
reg x_reg_23__retimed_I6442_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6442_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[8];
	end
assign N11530 = x_reg_23__retimed_I6442_QOUT;
reg x_reg_23__retimed_I6441_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6441_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993;
	end
assign N11528 = x_reg_23__retimed_I6441_QOUT;
reg x_reg_23__retimed_I6436_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6436_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5];
	end
assign N11515 = x_reg_23__retimed_I6436_QOUT;
reg x_reg_20__retimed_I6418_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6418_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7511;
	end
assign N11464 = x_reg_20__retimed_I6418_QOUT;
reg x_reg_20__retimed_I6417_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6417_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7473;
	end
assign N11462 = x_reg_20__retimed_I6417_QOUT;
reg x_reg_14__retimed_I6401_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6401_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490;
	end
assign N11418 = x_reg_14__retimed_I6401_QOUT;
reg x_reg_9__retimed_I6395_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I6395_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7467;
	end
assign N11401 = x_reg_9__retimed_I6395_QOUT;
reg x_reg_9__retimed_I6394_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I6394_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7433;
	end
assign N11399 = x_reg_9__retimed_I6394_QOUT;
reg x_reg_20__retimed_I6387_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6387_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7540;
	end
assign N11377 = x_reg_20__retimed_I6387_QOUT;
reg x_reg_21__retimed_I6385_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6385_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513;
	end
assign N11372 = x_reg_21__retimed_I6385_QOUT;
reg x_reg_21__retimed_I6383_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6383_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7493;
	end
assign N11368 = x_reg_21__retimed_I6383_QOUT;
reg x_reg_23__retimed_I6380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6380_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8206;
	end
assign N11360 = x_reg_23__retimed_I6380_QOUT;
reg x_reg_10__retimed_I6358_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I6358_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443;
	end
assign N11304 = x_reg_10__retimed_I6358_QOUT;
reg x_reg_17__retimed_I6356_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6356_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7532;
	end
assign N11299 = x_reg_17__retimed_I6356_QOUT;
reg x_reg_17__retimed_I6355_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6355_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7499;
	end
assign N11297 = x_reg_17__retimed_I6355_QOUT;
reg x_reg_17__retimed_I6353_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6353_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546;
	end
assign N11293 = x_reg_17__retimed_I6353_QOUT;
reg x_reg_19__retimed_I6352_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6352_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7517;
	end
assign N11290 = x_reg_19__retimed_I6352_QOUT;
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6824 (.Y(N12417), .A(N11290));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6825 (.Y(N12418), .A(N12417));
reg x_reg_19__retimed_I6351_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6351_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7479;
	end
assign N11288 = x_reg_19__retimed_I6351_QOUT;
reg x_reg_22__retimed_I6339_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6339_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7522;
	end
assign N11261 = x_reg_22__retimed_I6339_QOUT;
reg x_reg_2__retimed_I6300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I6300_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7481;
	end
assign N11143 = x_reg_2__retimed_I6300_QOUT;
reg x_reg_23__retimed_I6283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6283_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0];
	end
assign N11100 = x_reg_23__retimed_I6283_QOUT;
reg x_reg_22__retimed_I6275_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6275_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[46];
	end
assign N11079 = x_reg_22__retimed_I6275_QOUT;
reg x_reg_19__retimed_I6272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6272_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43];
	end
assign N11072 = x_reg_19__retimed_I6272_QOUT;
reg x_reg_18__retimed_I6269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I6269_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42];
	end
assign N11065 = x_reg_18__retimed_I6269_QOUT;
reg x_reg_17__retimed_I6266_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6266_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41];
	end
assign N11058 = x_reg_17__retimed_I6266_QOUT;
reg x_reg_15__retimed_I6263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I6263_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39];
	end
assign N11051 = x_reg_15__retimed_I6263_QOUT;
reg x_reg_14__retimed_I6260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6260_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38];
	end
assign N11044 = x_reg_14__retimed_I6260_QOUT;
reg x_reg_13__retimed_I6257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I6257_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37];
	end
assign N11037 = x_reg_13__retimed_I6257_QOUT;
reg x_reg_12__retimed_I6254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I6254_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36];
	end
assign N11030 = x_reg_12__retimed_I6254_QOUT;
reg x_reg_11__retimed_I6251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6251_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35];
	end
assign N11023 = x_reg_11__retimed_I6251_QOUT;
reg x_reg_9__retimed_I6248_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I6248_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33];
	end
assign N11016 = x_reg_9__retimed_I6248_QOUT;
reg x_reg_8__retimed_I6245_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I6245_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32];
	end
assign N11009 = x_reg_8__retimed_I6245_QOUT;
reg x_reg_5__retimed_I6242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I6242_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29];
	end
assign N11002 = x_reg_5__retimed_I6242_QOUT;
reg x_reg_4__retimed_I6239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I6239_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28];
	end
assign N10995 = x_reg_4__retimed_I6239_QOUT;
reg x_reg_0__retimed_I6236_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I6236_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24];
	end
assign N10988 = x_reg_0__retimed_I6236_QOUT;
reg x_reg_0__retimed_I6235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I6235_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[0];
	end
assign N10986 = x_reg_0__retimed_I6235_QOUT;
reg x_reg_21__retimed_I6233_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6233_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[45];
	end
assign N10981 = x_reg_21__retimed_I6233_QOUT;
reg x_reg_20__retimed_I6231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6231_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[44];
	end
assign N10976 = x_reg_20__retimed_I6231_QOUT;
reg x_reg_16__retimed_I6229_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I6229_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40];
	end
assign N10971 = x_reg_16__retimed_I6229_QOUT;
reg x_reg_10__retimed_I6227_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I6227_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34];
	end
assign N10966 = x_reg_10__retimed_I6227_QOUT;
reg x_reg_7__retimed_I6225_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I6225_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31];
	end
assign N10961 = x_reg_7__retimed_I6225_QOUT;
reg x_reg_6__retimed_I6223_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I6223_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30];
	end
assign N10956 = x_reg_6__retimed_I6223_QOUT;
reg x_reg_3__retimed_I6221_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I6221_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27];
	end
assign N10951 = x_reg_3__retimed_I6221_QOUT;
reg x_reg_2__retimed_I6219_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I6219_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26];
	end
assign N10946 = x_reg_2__retimed_I6219_QOUT;
reg x_reg_1__retimed_I6217_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I6217_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25];
	end
assign N10941 = x_reg_1__retimed_I6217_QOUT;
reg x_reg_23__retimed_I6213_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6213_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22678;
	end
assign N10901 = x_reg_23__retimed_I6213_QOUT;
reg x_reg_29__retimed_I6192_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__retimed_I6192_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8288;
	end
assign N10852 = x_reg_29__retimed_I6192_QOUT;
reg x_reg_0__retimed_I6186_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I6186_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8337;
	end
assign N10838 = x_reg_0__retimed_I6186_QOUT;
reg x_reg_1__retimed_I6183_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I6183_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8388;
	end
assign N10831 = x_reg_1__retimed_I6183_QOUT;
reg x_reg_2__retimed_I6180_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I6180_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8439;
	end
assign N10824 = x_reg_2__retimed_I6180_QOUT;
reg x_reg_3__retimed_I6177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I6177_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8483;
	end
assign N10817 = x_reg_3__retimed_I6177_QOUT;
reg x_reg_4__retimed_I6174_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I6174_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8533;
	end
assign N10810 = x_reg_4__retimed_I6174_QOUT;
reg x_reg_5__retimed_I6171_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I6171_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8360;
	end
assign N10803 = x_reg_5__retimed_I6171_QOUT;
reg x_reg_6__retimed_I6168_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I6168_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8408;
	end
assign N10796 = x_reg_6__retimed_I6168_QOUT;
reg x_reg_7__retimed_I6165_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I6165_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8457;
	end
assign N10789 = x_reg_7__retimed_I6165_QOUT;
reg x_reg_8__retimed_I6162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I6162_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8504;
	end
assign N10782 = x_reg_8__retimed_I6162_QOUT;
reg x_reg_9__retimed_I6159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I6159_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8553;
	end
assign N10775 = x_reg_9__retimed_I6159_QOUT;
reg x_reg_10__retimed_I6156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I6156_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8381;
	end
assign N10768 = x_reg_10__retimed_I6156_QOUT;
reg x_reg_11__retimed_I6153_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6153_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8429;
	end
assign N10761 = x_reg_11__retimed_I6153_QOUT;
reg x_reg_12__retimed_I6150_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I6150_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8474;
	end
assign N10754 = x_reg_12__retimed_I6150_QOUT;
reg x_reg_13__retimed_I6147_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I6147_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8522;
	end
assign N10747 = x_reg_13__retimed_I6147_QOUT;
reg x_reg_14__retimed_I6144_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6144_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8351;
	end
assign N10740 = x_reg_14__retimed_I6144_QOUT;
reg x_reg_15__retimed_I6141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I6141_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8400;
	end
assign N10733 = x_reg_15__retimed_I6141_QOUT;
reg x_reg_16__retimed_I6138_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I6138_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8450;
	end
assign N10726 = x_reg_16__retimed_I6138_QOUT;
reg x_reg_17__retimed_I6135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6135_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8494;
	end
assign N10719 = x_reg_17__retimed_I6135_QOUT;
reg x_reg_18__retimed_I6132_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I6132_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8543;
	end
assign N10712 = x_reg_18__retimed_I6132_QOUT;
reg x_reg_19__retimed_I6129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6129_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8371;
	end
assign N10705 = x_reg_19__retimed_I6129_QOUT;
reg x_reg_20__retimed_I6126_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6126_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8420;
	end
assign N10698 = x_reg_20__retimed_I6126_QOUT;
reg x_reg_21__retimed_I6123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6123_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8467;
	end
assign N10691 = x_reg_21__retimed_I6123_QOUT;
INVX3 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I0 (.Y(bdw_enable), .A(astall));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .A(b_man[19]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4362), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I3 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666), .A(a_man[19]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I4 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4063), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I5 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .A(b_man[20]));
CLKINVX4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144), .A(a_man[22]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I7 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3187), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I8 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3557), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3106), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4362), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4063), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3187));
INVX3 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I9 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .A(b_man[22]));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I10 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672), .A(a_man[21]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I11 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3808), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I12 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4090), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I13 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133), .A(a_man[20]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I14 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4967), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
CLKINVX4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I15 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .A(b_man[21]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I16 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4984), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I17 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5097), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4643), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4967), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4984));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I18 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3932), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3483), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3557), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3808), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4643));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I19 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4977), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I20 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4081), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I21 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .A(b_man[18]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I22 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4635), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6907 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184), .A(a_man[18]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I24 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3157), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I25 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3464), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I26 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3181), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4795), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4635), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3157), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3464));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I27 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4461), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4010), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4977), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4081), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3181));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I28 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3178), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I29 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4351), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I30 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4072), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I31 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4084), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3635), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3178), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4351), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4072));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I32 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3453), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I33 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4626), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I34 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4340), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I35 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4876), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4427), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3453), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4626), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4340));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I36 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .A(b_man[17]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I37 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4909), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I38 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715), .A(a_man[17]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I39 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4326), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I40 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3735), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I41 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3976), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3526), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4909), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4326), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3735));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I42 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4991), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4538), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4876), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3976), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4795));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I43 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3285), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4912), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3106), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4084), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4991));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I44 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3483), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4461), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3285));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I45 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .A(b_man[16]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I46 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3116), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I47 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176), .A(a_man[16]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I48 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3425), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I49 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4012), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I50 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3862), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3412), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3116), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3425), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4012));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I51 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3165), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I52 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3727), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I53 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4901), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I54 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4618), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I55 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4763), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4313), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3727), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4901), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4618));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I56 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3712), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3256), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3165), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4763));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I57 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4332), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I58 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3443), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I59 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .A(b_man[15]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I60 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3387), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I61 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .A(a_man[15]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I62 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4590), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I63 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4278), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I64 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4920), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4469), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3387), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4590), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4278));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I65 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3599), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3147), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4332), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3443), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4920));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I66 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4611), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4158), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4427), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3526), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3599));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I67 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3822), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3364), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3712), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3635), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4611));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I68 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3822), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4010), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4912));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I69 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I70 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4607), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I71 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3716), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I72 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3433), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I73 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4653), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4201), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4607), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3716), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3433));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I74 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4001), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I75 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3103), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I76 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4893), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I77 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3755), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3295), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4001), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3103), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4893));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I78 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4503), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4054), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3755), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3412));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I79 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4267), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I80 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3375), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I81 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3094), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I82 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3903), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3456), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4267), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3375), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3094));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I83 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .A(b_man[14]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I84 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3662), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I85 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232), .A(a_man[14]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I86 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3689), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I87 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4557), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I88 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5074), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4620), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3662), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3689), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4557));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I89 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4883), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I90 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3992), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I91 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3707), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I92 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4806), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4356), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4883), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3992), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3707));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I93 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3493), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5105), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3903), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5074), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4806));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I94 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3332), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4952), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3493), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4313), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3147));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I95 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3446), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5066), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3256), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4503), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3332));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I96 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4538), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3364));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I97 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I98 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I99 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4393), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3940), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3295), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4469), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4201));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I100 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3085), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I101 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4258), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I102 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3983), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I103 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4060), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3610), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3085), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4258), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3983));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I104 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4547), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4095), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4060), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3456));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I105 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .A(b_man[13]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I106 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3935), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I107 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758), .A(a_man[13]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I108 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4854), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I109 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4824), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I110 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4321), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3872), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3935), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4854), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4824));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I111 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4598), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I112 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4549), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I113 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3651), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I114 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3366), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I115 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3156), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4772), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4549), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3651), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3366));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I116 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3643), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3189), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4321), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4598), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3156));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I117 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3225), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4841), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4547), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3643), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5105));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I118 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4236), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3790), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4054), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4393), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3225));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I119 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4236), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4158), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5066));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I120 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I121 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3697), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I122 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4873), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I123 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .A(b_man[12]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I124 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4203), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I125 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220), .A(a_man[12]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I126 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3951), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I127 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5099), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I128 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4739), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4289), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4203), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3951), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5099));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I129 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4962), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4513), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3697), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4873), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4739));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I130 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3356), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I131 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I132 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4250), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I133 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4480), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4030), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3356), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4536), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4250));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I134 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4814), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I135 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3926), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I136 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3641), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I137 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3574), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3122), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4814), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3926), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3641));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I138 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3971), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I139 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5144), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I140 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4864), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I141 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3306), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4929), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3971), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5144), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4864));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I142 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3800), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3341), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4480), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3574), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3306));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I143 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3377), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4998), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4962), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4356), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3800));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I144 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4696), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4245), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4772), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3872), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3610));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I145 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4280), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3830), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4696), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3189), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4095));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I146 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4128), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3678), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3940), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3377), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4280));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I147 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4128), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4952), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3790));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I148 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I149 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I150 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I151 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5089), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I152 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4196), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I153 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3915), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I154 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3088), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4703), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5089), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4196), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3915));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I155 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .A(b_man[11]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I156 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4484), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I157 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .A(a_man[11]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I158 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5116), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I159 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3298), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I160 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4253), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3806), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4484), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5116), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3298));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I161 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3634), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I162 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4805), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I163 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4526), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I164 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3994), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3542), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3634), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4805), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4526));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I165 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4209), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3764), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3088), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4253), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3994));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I166 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4243), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I167 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3348), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I168 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5135), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I169 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4896), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3348), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5135));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I170 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5112), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4663), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4289), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4896), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3122));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I171 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3534), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3081), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4209), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5112));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I172 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .A(b_man[10]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I173 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4751), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I174 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273), .A(a_man[10]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I175 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4213), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I176 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3576), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I177 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4939), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4489), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4213), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3576));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I178 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3961), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I179 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4183), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I180 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4476), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I181 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3290), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I182 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3775), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3316), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4476), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4183), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3290));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I183 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3730), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3271), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4939), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3961), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3775));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I184 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3950), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3503), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4929), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4030), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3730));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I185 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4439), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3986), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3950), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3341), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4245));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I186 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3114), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4728), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4998), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3534), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4439));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I187 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3114), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4841), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3678));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I188 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I189 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3467), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5082), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3542), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4703), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4446));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I190 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4518), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I191 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3626), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I192 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3340), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I193 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3512), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5121), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4518), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3626), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3340));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I194 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3905), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I195 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5081), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I196 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4797), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I197 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4673), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4219), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3905), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5081), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4797));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I198 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4628), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4176), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3512), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4673), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3806));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I199 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4849), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4403), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3467), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4628), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3764));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I200 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5071), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I201 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3282), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I202 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4175), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I203 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4455), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4004), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5071), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3282), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4175));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I204 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4741), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I205 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3569), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I206 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4464), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I207 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3550), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3098), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4741), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3569), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4464));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I208 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4787), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I209 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3893), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I210 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3617), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I211 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3280), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4904), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4787), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3893), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3617));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I212 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3241), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4860), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4455), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3550), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3280));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I213 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5125), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I214 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4234), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I215 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .A(b_man[9]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I216 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5029), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I217 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801), .A(a_man[9]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I218 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3307), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I219 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3852), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I220 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4712), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4262), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5029), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3307), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3852));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I221 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4410), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3960), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5125), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4234), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4712));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I222 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3326), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I223 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4508), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I224 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4222), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I225 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4186), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3740), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3326), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4508), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4222));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I226 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4142), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3692), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4489), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4186), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3316));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I227 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4366), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3913), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3241), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4410), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4142));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I228 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3685), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3234), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4663), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4366));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I229 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3264), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4884), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3081), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4849), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3685));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I230 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3264), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3830), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4728));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I231 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I232 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I233 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3843), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I234 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5019), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I235 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4731), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I236 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4499), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4047), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5019), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3843), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4731));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I237 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .A(b_man[8]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I238 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3231), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I239 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260), .A(a_man[8]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I240 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4483), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I241 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4125), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I242 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3593), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3140), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3231), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4483), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4125));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I243 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4453), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I244 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3559), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I245 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3273), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I246 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3324), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4948), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3273), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3559), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4453));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I247 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5090), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4637), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4499), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3593), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3324));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I248 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5049), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4597), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5121), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4219), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5090));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I249 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3197), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4816), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4176), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3271), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5049));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I250 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3608), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I251 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4779), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I252 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4501), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I253 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5133), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4681), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3608), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4779), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4501));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I254 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5065), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I255 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4169), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I256 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3885), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I257 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4229), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3784), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5065), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4169), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3885));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I258 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3924), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3476), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5133), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4229), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4262));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I259 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4826), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4376), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4004), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4904), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3098));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I260 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3881), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3428), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3960), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3924), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4826));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I261 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4103), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3653), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3881), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5082), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3913));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I262 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4589), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4135), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4403), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3197), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4103));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I263 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4589), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3986), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4884));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I264 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I265 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .A(b_man[7]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I266 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3508), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I267 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792), .A(a_man[7]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I268 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3579), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I269 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4400), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I270 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3638), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3184), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3508), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3579), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4400));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I271 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3317), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I272 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5009), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I273 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4114), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I274 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3223), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I275 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4543), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4086), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5009), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4114), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3223));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I276 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3969), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3521), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3638), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3317), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4543));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I277 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3263), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I278 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4160), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I279 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4445), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I280 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4274), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3825), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3263), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4160), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4445));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I281 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4724), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I282 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3832), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I283 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3549), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I284 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3368), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4994), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4724), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3832), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3549));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I285 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3876), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I286 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5055), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I287 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4770), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I288 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3110), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4722), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3876), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5055), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4770));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I289 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4869), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4420), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4274), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3368), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3110));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I290 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3664), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3207), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3969), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3740), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4869));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I291 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4780), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4328), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3692), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4860), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3664));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I292 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3705), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3250), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4948), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3140), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4047));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I293 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4493), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I294 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3597), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I295 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .A(b_man[6]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I296 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3781), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I297 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318), .A(a_man[6]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I298 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4740), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I299 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4668), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I300 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4843), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4397), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3781), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4740), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4668));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I301 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4014), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3561), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4493), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3597), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4843));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I302 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4605), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4153), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4681), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3784), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4014));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I303 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4564), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4112), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4637), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3705), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4605));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I304 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3621), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3163), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4564), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4597), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3428));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I305 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5006), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4555), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4816), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4780), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3621));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I306 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5006), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3234), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4135));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I307 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I308 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I309 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I310 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4760), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I311 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3869), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I312 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3587), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I313 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3150), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4767), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4760), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3869), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3587));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I314 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4150), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I315 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3254), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I316 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5047), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I317 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4316), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3867), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4150), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3254), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5047));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I318 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3749), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3288), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3150), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4316), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I319 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5001), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I320 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4105), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I321 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3824), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I322 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4581), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4131), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4105), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5001), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3824));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I323 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4389), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I324 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3501), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I325 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3212), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I326 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3681), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3228), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3501), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4389), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3212));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I327 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4714), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I328 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3541), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I329 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4436), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I330 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3415), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5036), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4436), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3541), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4714));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I331 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4915), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4465), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4581), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3681), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3415));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I332 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3439), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5059), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3749), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4915), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3521));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I333 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3397), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5017), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3476), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3439));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I334 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4646), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4197), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4994), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4086), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3825));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I335 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4339), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3889), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4420), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4646), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3250));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I336 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4299), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3848), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4339), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3207), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4112));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I337 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4520), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4067), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4328), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3397), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I338 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4520), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3653), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4555));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I339 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I340 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .A(b_man[5]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I341 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4052), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I342 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845), .A(a_man[5]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I343 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3842), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I344 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4942), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I345 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3084), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4699), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4052), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3842), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4942));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I346 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4098), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I347 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3202), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I348 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4378), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I349 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4888), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4098), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3202), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4378));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I350 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4660), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I351 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3774), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I352 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3490), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I353 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3990), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3537), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3774), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3490));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I354 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4056), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3602), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3084), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4888), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3990));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I355 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3245), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I356 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I357 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4426), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I358 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4623), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4170), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3245), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4426), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3536));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I359 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3814), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I360 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4993), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I361 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4705), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I362 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3726), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3267), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3814), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4993), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4705));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I363 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5039), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I364 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4141), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I365 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3859), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I366 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3459), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5078), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5039), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4141), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3859));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I367 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4956), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4507), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4623), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3726), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3459));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I368 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3488), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5100), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4056), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4722), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4956));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I369 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3793), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3337), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4397), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4131));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I370 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4386), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3933), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3793), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3561), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4465));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I371 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3174), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4789), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4153), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3488), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4386));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I372 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4690), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4239), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3867), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4767), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5036));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I373 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3217), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4835), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4690), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3288), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4197));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I374 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4077), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3628), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5059), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3889));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I375 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3131), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4749), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5017), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3174), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4077));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I376 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3163), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4067));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I377 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I378 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I379 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5003), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4551), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4170), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4442), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3267));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I380 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4431), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3980), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3602), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5003), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4507));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I381 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4982), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I382 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3191), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I383 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4088), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I384 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3125), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4743), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4982), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3191), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4088));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I385 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3528), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I386 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4695), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I387 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3805), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I388 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4033), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3578), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3528), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4695), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3805));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I389 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4368), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I390 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3478), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I391 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4650), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I392 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4294), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3841), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3478), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4650));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I393 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3193), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4808), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3125), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4033), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4294));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I394 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4750), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I395 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4043), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I396 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4935), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I397 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3760), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I398 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3392), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5011), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4043), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4935), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3760));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I399 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299), .A(a_man[4]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I400 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5012), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I401 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3146), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I402 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737), .A(b_man[4]));
CLKINVX4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I403 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11793), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I404 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11793));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I405 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4320), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I406 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4559), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4107), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5012), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3146), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4320));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I407 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4361), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3909), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4750), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3392), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4559));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I408 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3238), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I409 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4417), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I410 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4133), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I411 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4934), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4482), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3238), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4417), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4133));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I412 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4096), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3647), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4934), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4699), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3537));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I413 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3529), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5143), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3193), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4361), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4096));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I414 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4123), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3673), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4431), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3529), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5100));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I415 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3851), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I416 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5031), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I417 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835), .A(a_man[3]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I418 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4104), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
CLKINVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I419 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .A(b_man[3]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I420 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4596), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I421 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3420), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I422 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5124), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4675), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4104), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4596), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3420));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I423 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3768), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3309), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5031), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5124));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I424 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4927), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I425 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3752), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I426 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4640), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I427 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4863), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4413), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4927), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3752), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4640));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I428 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3138), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I429 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4312), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I430 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4036), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I431 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3963), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3515), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3138), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4312), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4036));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I432 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4359), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I433 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3183), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I434 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3469), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I435 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3696), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3244), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4359), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3183), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3469));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I436 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4666), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4212), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4863), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3963), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3696));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I437 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3833), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3379), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5078), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3768), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4666));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I438 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3258), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4878), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3833), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4239), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3337));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I439 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5027), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4572), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3933), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3258), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4835));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I440 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4983), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4532), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4123), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4789), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5027));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I441 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4983), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3848), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4749));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I442 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I443 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4685), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I444 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3519), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I445 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4409), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I446 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3432), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5051), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4685), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3519), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4409));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I447 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4079), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I448 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4973), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I449 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3797), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I450 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4600), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4147), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4079), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4973), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3797));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I451 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4124), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I452 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3230), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I453 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5021), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I454 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4331), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3884), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4124), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3230), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5021));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I455 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3507), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5115), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4600), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4331));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I456 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4729), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4284), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3909), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3507), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4808));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I457 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3237), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4853), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4743), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4482));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I458 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4406), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3953), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4107), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5011), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3841));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I459 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3570), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3118), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3237), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4406), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3647));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I460 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4161), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3715), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4729), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3570), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5143));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I461 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4348), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I462 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3172), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I463 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4069), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I464 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4265), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3817), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4348), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3172), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4069));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I465 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4633), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I466 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3742), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I467 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3461), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I468 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3361), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4986), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4633), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3742), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3461));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I469 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3789), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I470 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4964), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I471 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4676), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I472 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3101), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4716), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3789), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4964), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4676));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I473 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4071), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3622), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4265), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3361), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3101));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I474 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4026), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I475 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4916), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I476 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3130), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I477 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4535), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4080), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4026), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4916), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3130));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6908 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .A(b_man[2]));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I479 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4868), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811));
CLKINVX4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I480 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934), .A(a_man[2]));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I481 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3201), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I482 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3695), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I483 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4792), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4342), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4868), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3201), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3695));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I484 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3410), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I485 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4587), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I486 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4302), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I487 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3631), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3177), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3410), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4587), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4302));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I488 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3167), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4784), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4535), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4792), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3631));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I489 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4139), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3688), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4071), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3167), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3309));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I490 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4474), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4020), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4551), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4139), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3379));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I491 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5068), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4615), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4474), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3980), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4878));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I492 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3855), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3406), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3673), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4161), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5068));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I493 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3628), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3855), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4532));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I494 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I495 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I496 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I497 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866));
OR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I498 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3786), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I499 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4514), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I500 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3623), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I501 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3334), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I502 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5075), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4621), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4514), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3623), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3334));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I503 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5079), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I504 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4793), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I505 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3900), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I506 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4168), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3719), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5079), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4793), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3900));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I507 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5123), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I508 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4231), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
CLKINVX4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I509 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891), .A(a_man[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I510 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3946), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I511 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3904), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3457), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5123), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4231), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3946));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I512 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4502), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4055), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5075), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4168), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3904));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I513 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .A(b_man[0]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I514 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5042), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
CLKINVX8 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I515 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .A(b_man[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I516 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3865), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I517 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3494), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5106), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5042), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3865));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I518 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3874), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I519 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4766), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I520 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4344), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3896), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3874), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4766));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I521 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3582), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I522 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4757), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I523 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4479), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I524 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4394), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3937), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3582), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4757), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4479));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I525 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4462), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4011), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3494), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3896), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4394));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I526 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3629), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I527 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3911), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I528 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4803), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I529 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4129), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3679), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3629), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3911), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4803));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I530 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4190), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I531 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5087), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I532 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3294), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I533 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3224), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4842), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4190), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5087), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3294));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I534 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3333), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4953), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3679), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4842), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3937));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I535 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4833), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4383), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4502), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4011), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3333));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I536 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3287), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I537 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4468), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I538 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4181), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I539 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3265), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4885), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3287), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4468), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4181));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I540 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3374), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4999), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3719), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4621), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4885));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I541 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4748), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I542 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3857), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I543 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3573), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I544 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4435), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3987), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4748), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3857), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3573));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I545 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3600), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3144), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5106), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4435), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3265));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I546 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3977), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3527), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4055), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3374), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3144));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I547 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4165), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I548 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3269), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I549 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5061), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I550 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4894), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4447), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4165), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3269), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5061));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I551 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4451), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I552 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4727), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I553 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3554), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I554 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3995), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3540), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4451), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4727), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3554));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I555 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4774), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I556 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3882), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I557 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3604), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I558 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3731), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3272), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4774), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3882), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3604));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I559 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4585), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4136), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4894), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3995), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3731));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I560 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3235), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I561 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4130), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I562 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4481), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4028), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3235), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4130));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I563 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4405), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I564 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3227), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I565 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4251), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3807), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4405), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3227));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I566 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5016), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I567 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4122), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I568 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3838), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I569 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3089), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4704), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5016), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4122), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3838));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I570 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3686), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3232), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4028), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4251), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3089));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I571 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4281), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3831), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4585), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3457), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3686));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I572 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3957), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I573 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5131), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I574 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4847), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I575 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3860), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3413), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3957), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5131), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4847));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I576 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3343), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I577 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4522), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I578 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4241), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I579 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5034), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4575), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3343), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4522), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4241));
CLKINVX4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I580 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346), .A(a_man[0]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I581 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4838), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I582 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4138), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I583 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5035), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I584 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3535), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3079), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4138), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5035));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I585 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4804), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4357), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4838), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4481), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3079));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I586 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4237), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3788), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3413), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4575), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4804));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I587 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4877), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4425), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4953), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4281), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3788));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I588 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3403), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5024), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4383), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3977), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4877));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I589 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3873), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I590 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5052), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I591 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4765), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I592 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4411), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3956), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3873), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5052), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4765));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I593 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3261), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I594 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4443), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I595 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4156), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I596 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3513), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5122), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3261), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4443), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4156));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I597 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4367), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3914), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4411), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3513), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I598 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3216), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I599 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4111), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I600 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5005), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I601 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3776), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3312), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3216), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4111), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5005));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I602 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4718), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I603 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3829), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I604 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3547), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I605 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4671), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4220), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4718), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3829), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3547));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I606 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3465), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5083), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3807), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3776), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4671));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I607 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3198), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4813), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3540), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3272));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I608 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3153), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4773), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4367), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3465), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3198));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I609 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3313), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I610 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4497), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I611 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3505), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I612 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4396), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I613 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4940), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4490), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3505), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4396));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I614 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4629), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4174), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3313), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4497), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4940));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I615 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3847), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I616 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5026), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I617 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4736), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I618 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3302), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4930), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3847), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5026), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4736));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I619 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4458), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I620 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3563), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I621 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3277), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I622 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4210), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3765), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4458), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3563), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3277));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I623 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3422), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5041), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4629), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4930), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3765));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I624 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4061), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3611), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3232), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4136), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5041));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I625 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4921), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4470), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3831), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3153), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4061));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I626 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4612), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4159), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4425), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3527), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4921));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I627 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3286), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4908), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3224), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4129), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5034));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I628 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4488), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I629 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3303), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I630 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3592), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I631 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3182), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4796), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4488), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3303), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3592));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I632 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4569), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I633 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3680), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I634 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4764), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4314), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4569), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3680), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3535));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I635 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4194), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3747), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3860), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4796), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4764));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I636 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3671), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3214), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4237), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4908), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3747));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I637 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5069), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I638 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4173), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I639 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3891), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I640 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5113), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4661), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5069), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4173), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3891));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I641 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3644), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3190), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5113), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3302), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4210));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I642 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3614), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I643 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4782), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I644 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4505), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I645 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3945), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3504), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3614), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4782), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4505));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I646 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4216), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I647 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3322), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I648 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5114), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I649 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4850), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4404), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4216), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3322), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5114));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I650 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4548), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4093), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3945), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4850), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3987));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I651 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5138), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4689), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3644), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4314), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4548));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I652 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4811), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I653 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3639), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I654 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4534), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I655 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4988), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4539), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3639), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4534));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I656 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5094), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I657 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4199), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I658 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3920), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I659 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4085), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3633), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5094), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4199), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3920));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I660 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4248), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I661 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5141), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I662 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3352), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I663 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3823), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3365), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4248), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5141), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3352));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I664 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5098), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4644), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4539), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3633), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3365));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I665 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3399), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I666 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4576), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I667 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4295), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I668 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3553), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3107), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4576), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4295));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I669 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4858), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I670 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3687), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I671 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3967), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I672 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4721), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4266), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3687), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4858), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3967));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I673 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3929), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3484), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3107), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4266), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3600));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I674 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4568), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4120), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5138), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4644), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3484));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I675 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3115), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4726), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3422), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4357), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3190));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I676 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4322), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3870), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4661), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4404));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I677 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4018), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3566), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4322), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4093), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4999));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I678 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3710), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3257), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4689), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3115), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4018));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I679 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4304), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3853), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3214), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4120), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3710));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I680 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5024), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4612), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3853));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I681 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3888), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3437), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4721), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3823), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3553));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I682 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5054), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4603), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4085), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3182), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4988));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I683 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3355), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4979), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3437), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4603), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4194));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I684 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4000), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3546), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4979), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3671), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4568));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I685 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3082), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I686 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3979), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I687 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4255), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I688 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3518), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5127), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3082), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3979), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4255));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I689 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3694), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I690 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4871), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I691 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4586), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I692 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4416), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3966), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4586), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4871), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3694));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I693 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4305), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I694 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3409), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I695 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3129), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I696 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3248), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4866), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4305), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3409), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3129));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I697 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3625), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3171), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5127), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3966), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4866));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I698 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4025), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I699 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3601), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I700 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4775), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
ADDHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I701 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4046), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3590), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3601), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4775));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I702 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4149), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3699), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4344), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4025), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3590));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I703 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4529), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4074), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3286), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4462), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3699));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I704 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3096), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4710), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4833), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3171), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4074));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I705 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3314), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6909 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4498), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I707 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4208), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I708 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4944), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4494), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3314), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4498), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4208));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I709 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3930), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I710 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5104), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I711 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4822), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I712 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3779), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3321), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3930), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5104), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4822));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I713 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4545), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I714 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3649), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I715 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3362), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I716 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4679), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4225), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4545), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3649), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3362));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I717 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4786), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4334), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4494), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3321), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4225));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I718 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4257), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3813), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3929), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5098), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4334));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I719 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4900), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4452), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4710), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3813), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3403));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I720 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3546), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4304), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4452));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I721 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I722 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4487), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4034), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4679), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3518), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4416));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I723 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3612), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I724 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4506), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I725 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4634), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4180), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3612), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4506));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I726 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3581), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3128), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4180), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4944), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3779));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I727 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4856), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4408), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4034), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3625), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3128));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I728 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4553), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I729 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3372), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I730 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4263), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I731 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3205), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4821), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4553), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3372), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4263));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I732 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3988), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I733 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3091), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I734 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4880), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I735 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4109), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3661), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3091), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4880));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I736 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4595), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I737 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3703), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I738 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3419), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I739 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5014), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4563), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4595), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3703), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3419));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I740 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4215), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3772), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4821), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3661), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4563));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I741 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4217), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I742 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3323), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I743 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5111), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I744 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3472), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5088), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3323), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5111));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I745 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3659), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I746 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3938), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I747 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4829), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I748 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4373), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3922), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3659), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4829), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3938));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I749 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3311), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4937), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3248), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5088), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3922));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I750 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3691), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3239), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3772), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4937), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4529));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I751 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3426), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5046), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4408), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4257), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3239));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I752 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3137), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I753 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4315), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I754 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4035), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I755 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3846), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3393), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3137), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4315), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4035));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I756 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5119), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4670), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4149), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3393), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5054));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I757 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4926), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I758 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3754), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I759 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4744), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4298), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4926), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3754), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4046));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I760 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3955), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3510), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4298), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3888), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4786));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I761 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4592), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4140), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3355), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4670), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3510));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I762 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4327), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3877), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4140), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3096), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4000));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I763 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4900), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5046), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3877));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I764 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743));
AND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I765 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I766 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3947), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I767 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4228), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I768 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5120), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I769 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4969), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4519), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3947), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5120));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I770 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4810), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4363), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3846), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5014), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4519));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I771 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4839), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I772 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3668), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I773 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4561), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704));
ADDFHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I774 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3804), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3347), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4839), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3668), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4561));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I775 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4275), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I776 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3100), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I777 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3384), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I778 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4702), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4249), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3100), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4275), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3384));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I779 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3650), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3195), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3347), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4249), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4744));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I780 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3121), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4733), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4363), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4215), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3195));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I781 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3761), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3300), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4733), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3691), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4592));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I782 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4649), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I783 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3762), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I784 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3477), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I785 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4172), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3728), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4649), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3762), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3477));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I786 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3383), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5004), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3581), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3728), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4487));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I787 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3912), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3463), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4109), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3205), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4373));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I788 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4515), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I789 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3335), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I790 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4065), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3616), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4515), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3335));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I791 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5080), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4625), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4634), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3472));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I792 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4287), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3836), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4625), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3311));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I793 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4928), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4478), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5004), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4856), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3836));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I794 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3430), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I795 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4323), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I796 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4604), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I797 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4444), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3991), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4323), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3430), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4604));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I798 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4890), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I799 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3996), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I800 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3714), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I801 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3538), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3086), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4890), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3996), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3714));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I802 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4042), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I803 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4938), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I804 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3145), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I805 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3270), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4892), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4042), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4938), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3145));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I806 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4554), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4099), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3991), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3086), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4892));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I807 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4024), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3571), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4099), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5119), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3955));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I808 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4658), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4207), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4478), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3571), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3426));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I809 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4327), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3300), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4207));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I810 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I811 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3344), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I812 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5132), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I813 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3958), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I814 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3229), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4846), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3344), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5132), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3958));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I815 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4570), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I816 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3677), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I817 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4848), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I818 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4134), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3683), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4570), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3677), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4848));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I819 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3982), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3532), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4846), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4172), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3683));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I820 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4898), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I821 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4008), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I822 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3724), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I823 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3868), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3417), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4898), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4008), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3724));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I824 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3112), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I825 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3394), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I826 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4285), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I827 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5038), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4582), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3394), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3112), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4285));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I828 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3441), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I829 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4613), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I830 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4330), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I831 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4769), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4319), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3441), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4613), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4330));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I832 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4882), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4433), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4582), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4319));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I833 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4352), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3901), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4554), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3532), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4433));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I834 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4659), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I835 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3773), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I836 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3489), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I837 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4510), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4058), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4659), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3773), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3489));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I838 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4051), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I839 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3154), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I840 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4945), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I841 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3607), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3152), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4051), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3154), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4945));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I842 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3717), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3262), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4058), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3152), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3912));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I843 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3186), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4802), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3383), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3262), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4287));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I844 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4995), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4546), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3901), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4024), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4802));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I845 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4380), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I846 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3468), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I847 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4238), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I848 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4401), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3944), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3468), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4238));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I849 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3339), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4959), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4065), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4380), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3944));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I850 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4617), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4164), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5080), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4810), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4959));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I851 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4242), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3795), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3804), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4702), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4969));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I852 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5145), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4693), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4444), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3270), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3538));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I853 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3452), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5070), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3650), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3795), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4693));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I854 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4089), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3640), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3121), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4164), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5070));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I855 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3828), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3370), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3640), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4928), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3761));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I856 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4658), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4546), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3370));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I857 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739));
CLKAND2X3 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I858 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759));
NAND2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I859 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22954), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I860 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4664), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I861 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3496), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I862 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4456), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4005), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4664), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3496));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I863 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3767), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I864 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4655), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I865 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4870), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4419), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3767), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4655));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I866 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4374), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I867 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3486), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I868 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3196), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I869 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3702), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3251), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4374), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3486), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3196));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I870 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4823), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4377), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4005), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4870), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3702));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I871 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3878), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3429), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3956), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5122), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4823));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I872 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3533), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I873 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4701), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I874 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4422), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I875 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3440), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5057), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3533), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4701), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4422));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I876 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4989), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I877 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4094), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I878 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3811), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I879 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4606), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4154), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4989), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4094), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3811));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I880 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3206), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I881 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4385), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I882 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4102), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I883 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3281), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4902), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3206), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4385), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4102));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I884 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3665), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3208), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3440), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4606), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4902));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I885 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3539), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I886 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3252), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I887 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4432), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I888 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5091), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4638), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3539), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3252), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4432));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I889 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4137), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I890 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3242), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I891 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3757), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I892 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4932), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I893 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4121), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3674), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3757), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4932));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I894 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4337), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3890), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4137), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3242), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4121));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I895 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3819), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I896 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11781), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I897 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4709), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I898 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4182), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3741), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3819), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11781), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4709));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I899 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4565), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4110), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4638), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4337), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3741));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I900 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4300), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3849), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4377), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3208), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4110));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I901 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3595), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I902 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3240), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4861), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4456), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3595), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4490));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I903 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4143), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3693), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5091), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4182), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3281));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I904 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4781), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4329), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3665), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3693));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I905 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4521), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4068), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3429), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4300), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4329));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I906 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4101), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3654), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4174), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3240), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4143));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I907 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3840), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3386), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3878), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4813), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3654));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I908 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5044), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I909 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4145), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I910 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3864), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I911 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3925), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3474), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5044), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4145), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3864));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I912 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5050), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4594), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3312), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3925), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4220));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I913 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5007), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4556), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5050), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5083), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3914));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I914 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4645), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I915 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3475), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I916 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4365), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I917 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5028), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4573), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4645), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3475), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4365));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I918 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4082), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I919 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3188), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I920 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4980), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I921 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3856), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3405), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4082), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3188), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4980));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I922 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3175), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4790), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5028), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4419), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3856));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I923 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4692), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I924 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3803), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I925 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3523), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I926 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4756), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4308), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4692), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3803), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3523));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I927 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4078), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3627), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4756), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3251), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4154));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I928 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3396), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5018), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3175), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3474), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4078));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I929 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3619), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3164), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4594), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4565), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3396));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I930 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4734), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4290), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4556), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4781), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3619));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I931 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4521), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3386), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4290));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I932 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4963), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4511), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4101), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3870), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5007));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I933 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3796), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3342), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4773), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3840));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I934 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4734), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4511), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3342));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I935 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I936 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3756), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3293), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4726), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4963));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I937 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3796), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4470), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3293));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I938 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I939 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I940 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3756), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3257), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4159));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I941 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I942 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I943 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I944 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22921), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I945 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3325), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4949), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3405), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4573));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I946 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3816), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3360), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3325), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3890), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4790));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I947 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4031), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I948 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4923), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I949 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4271), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3826), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4031), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4923));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I950 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4414), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I951 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3594), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3141), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4271), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4414), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3674));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I952 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3794), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I953 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4970), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I954 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4683), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I955 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4913), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4466), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4970), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4683));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I956 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3179), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I957 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4354), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I958 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4073), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I959 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4015), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3558), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3179), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4354), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4073));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I960 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4636), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I961 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3748), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I962 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3466), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I963 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3111), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4723), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4636), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3748), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3466));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I964 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4496), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4048), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4913), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4015), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3111));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I965 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4981), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4533), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3594), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5057), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4496));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I966 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3132), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4747), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3816), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4981), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5018));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I967 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3164), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3132), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4068));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I968 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I969 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3124), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I970 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4022), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I971 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3259), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4879), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3124), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4022));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I972 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4335), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I973 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4619), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I974 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3444), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I975 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4957), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4504), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4335), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3444), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4619));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I976 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4903), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I977 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4013), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I978 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3729), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I979 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4057), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3603), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4903), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4013), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3729));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I980 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4800), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4347), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4879), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4957), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4057));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I981 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3485), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5101), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4466), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3558), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4800));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I982 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4345), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I983 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3458), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I984 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3168), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I985 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5067), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4616), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4345), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3458), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3168));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I986 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4960), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I987 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4064), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I988 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4292), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I989 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3117), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I990 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3148), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4768), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4292), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3117));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I991 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3899), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3450), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4960), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4064), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3148));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I992 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4647), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4195), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5067), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3899), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4723));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I993 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5130), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4682), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3485), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4647), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4949));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I994 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3738), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I995 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4914), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I996 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4627), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I997 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4162), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3713), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3738), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4914), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4627));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I998 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3750), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3289), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3826), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3259), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4162));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I999 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4230), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3783), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3141), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3750), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4048));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1000 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4713), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4259), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3627), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4230));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1001 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5130), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3360), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4259));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1002 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3849), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4747));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1003 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1004 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1005 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22578), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1006 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3160), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1007 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3389), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1008 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4283), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1009 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3941), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3499), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3389), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4283));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1010 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3791), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3338), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3160), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3941), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4768));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1011 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3636), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3185), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3713), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3791));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1012 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4387), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3934), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3636), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3289), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4195));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1013 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3783), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4387), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4682));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1014 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1015 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4609), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1016 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3720), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1017 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3435), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1018 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3682), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3226), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4609), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3720), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3435));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1019 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4003), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1020 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3108), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1021 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4895), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1022 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4844), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4398), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4003), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3108), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4895));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1023 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4691), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4240), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3682), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4844), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3603));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1024 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4544), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4087), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4691), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3450), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4347));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1025 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4544), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5101), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3934));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1026 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1027 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4558), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1028 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3378), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1029 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3568), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3119), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4558), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3378));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1030 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3097), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1031 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4272), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1032 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3993), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1033 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4475), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4021), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3097), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4272), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3993));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1034 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4579), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4132), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3499), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3568), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4475));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1035 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3530), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5140), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4579), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4504), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3338));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1036 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3185), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3530), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4087));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1037 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1038 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4477), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1039 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4260), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1040 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3367), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1041 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3087), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1042 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5000), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4552), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4260), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3367), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3087));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1043 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3358), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1044 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4541), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1045 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4252), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1046 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4358), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3910), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3358), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4541), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4252));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1047 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3917), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1048 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4807), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1049 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3723), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3917), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4807));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1050 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4817), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1051 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3646), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1052 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3460), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5076), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4817), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3646));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1053 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3194), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3723), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5076), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3910));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1054 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4552), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4358), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3194));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1055 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3711), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1056 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4886), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1057 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3656), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1058 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4550), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1059 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4097), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3645), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3656), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4550));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1060 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3297), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4925), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3711), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4886), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4097));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1061 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3985), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1062 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3834), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3460), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3985), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3645));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1063 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4206), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3759), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5000), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3119), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4021));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1064 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4925), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3834), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3759));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1065 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1066 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1067 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3700), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1068 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4531), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1069 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3637), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1070 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5084), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1071 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3907), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1072 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4889), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5084), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3907));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1073 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4531), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3637), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4889));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1074 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1075 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1076 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4680), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1077 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1078 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1079 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1080 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1081 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1082 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1083 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1084 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1085 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4226), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1086 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4680), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4226));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1087 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1088 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1089 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1090 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3249), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943));
OAI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1091 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3700), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3249));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1092 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1093 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1094 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3416), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5037), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3226), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4398), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3297));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1095 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4132), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4206), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5037));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1096 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1097 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4530), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1098 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1099 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4075), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678));
OAI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1100 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4530), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4075));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1101 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4240), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3416), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5140));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1102 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1103 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1104 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3737), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1105 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1106 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1107 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3279), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1108 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3279));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1109 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1110 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1111 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4027), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148));
OAI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1112 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4477), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4027));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1113 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1114 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1115 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1116 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1117 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22570), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566));
OAI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1118 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22578), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22570));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1119 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1120 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5045), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1121 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5045));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1122 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1123 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1124 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1125 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1126 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1127 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4516), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146));
OAI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1128 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22911), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4516));
AOI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1129 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22921), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22911));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1130 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1131 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1132 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22737), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1133 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22737));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1134 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1135 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1136 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22745), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1137 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22922), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22745));
AOI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1138 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22934), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22922));
OAI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1139 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22954), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22934));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1140 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4402), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1141 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11813), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1142 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3222), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1143 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4007), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3552), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4402), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11813), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3222));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1144 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4976), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4525), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4007), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3515), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4675));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1145 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3810), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3354), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4413), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3244), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4147));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1146 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5043), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4591), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4976), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3810));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1147 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4371), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1148 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3968), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1149 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3562), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3113), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4371), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3968));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1150 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4113), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1151 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5142), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1152 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3684), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1153 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4859), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1154 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4467), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4016), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5142), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3684), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4859));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1155 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4907), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4457), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3562), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4113), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4467));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1156 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4707), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4254), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3884), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5051), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4907));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1157 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3875), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3424), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4707), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5115), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3953));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1158 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3296), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4924), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5043), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3875), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4284));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1159 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4954), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1160 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3780), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1161 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4667), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1162 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4836), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4390), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4954), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3780), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4667));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1163 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4059), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1164 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3162), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1165 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4338), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1166 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3936), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3491), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4059), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3162), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4338));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1167 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4391), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1168 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3500), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1169 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3211), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1170 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3675), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3221), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3500), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3211));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1171 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4639), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4188), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4836), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3936), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3675));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1172 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4017), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1173 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3120), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1174 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4905), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1175 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4198), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3753), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4017), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3120), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4905));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1176 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4622), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1177 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3732), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1178 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3451), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1179 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5102), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4648), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4622), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3732), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3451));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1180 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4577), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1181 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3400), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1182 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4296), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1183 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3291), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4917), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4577), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3400), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4296));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1184 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3743), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3283), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4198), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5102), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3291));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1185 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3480), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5092), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4080), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4342), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3177));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1186 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3543), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3093), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4639), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3743), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3480));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1187 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4379), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3927), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3817), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4716), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4986));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1188 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4450), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3998), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4784), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3622), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4379));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1189 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4777), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4325), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3543), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4450));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1190 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4205), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3758), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4777), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3118), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4020));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1191 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3898), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3449), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3715), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3296), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4205));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1192 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3898), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4572), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3406));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1193 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1194 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4574), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4126), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3113), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4401), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3229));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1195 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3407), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5030), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5038), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4134), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3868));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1196 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3210), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4828), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4574), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3552), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3407));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1197 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3276), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4897), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3210), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4525), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3354));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1198 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3613), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3159), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4591), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3688), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3276));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1199 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4311), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3858), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3607), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4510), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4769));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1200 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3142), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4761), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3753), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4016), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4917));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1201 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4115), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3667), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4311), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4457), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3142));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1202 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4049), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3596), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4648), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4390), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3491));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1203 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5020), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4566), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4049), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3283), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4188));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1204 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4177), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3734), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4115), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4254), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5020));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1205 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4517), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4062), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3424), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4177), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4325));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1206 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5107), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4657), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3613), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4517));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1207 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5107), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4615), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3449));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1208 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307));
CLKAND2X3 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1209 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1210 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4950), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4500), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3339), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3221), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4242));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1211 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3850), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3398), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4950), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5092), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3927));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1212 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5086), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4632), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3093), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3850), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3998));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1213 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3785), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3327), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5145), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4126), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5030));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1214 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4684), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4233), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3982), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3858), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4882));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1215 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4752), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4301), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4828), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3785), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4684));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1216 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3918), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3471), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4897), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4752), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3734));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1217 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3345), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4966), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3159), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5086), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3918));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1218 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3345), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3758), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4657));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1219 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1220 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3524), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5134), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4761), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3717), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3596));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1221 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3586), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3134), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3667), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3524));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1222 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4421), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3972), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4617), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4500), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3452));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1223 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4492), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4041), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3398), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4421), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4301));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1224 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4819), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4370), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4632), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3586), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4492));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1225 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4819), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4062), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4966));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1226 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498));
CLKAND2X3 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1227 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449));
NAND2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1228 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1229 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4155), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3706), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3186), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3972));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1230 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3253), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4872), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4233), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3327), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4352));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1231 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5060), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4608), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4872), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4089), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4995));
ADDFXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1232 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3828), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3706), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4608));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1233 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1234 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3318), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4941), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3253), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4155));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1235 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5060), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4041), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4941));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1236 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777));
CLKAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1237 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809));
ADDFHXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1238 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3471), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4370));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1239 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1240 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200));
CLKAND2X3 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1241 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1242 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1243 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22928), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1244 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1245 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1246 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3192), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1247 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3192));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1248 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1249 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1250 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5002), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1251 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22938), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5002));
AOI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1252 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22938));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1253 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1254 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1255 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4732), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1256 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4732));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1257 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1258 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1259 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4473), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1260 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22919), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4473));
AOI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1261 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22947), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22919));
OAI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1262 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22917), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22947));
AOI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1263 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22928), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22917));
NOR2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1264 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1265 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1266 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1267 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1268 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1269 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3942), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106));
OAI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1270 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3942));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1271 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1272 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1273 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1274 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1275 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1276 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4958), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577));
OAI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1277 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4430), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4958));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1278 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4430));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1279 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1280 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1281 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1282 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1283 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1284 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3897), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117));
OA21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1285 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5032), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3897));
OAI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1286 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3427), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5032));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1287 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3328), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3427));
OAI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6899 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3786), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3328));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1289 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1290 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3818), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1291 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3801), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1292 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4708), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1293 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3670), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3215), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3818), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3801), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4708));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1294 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3215), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5097), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3932));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1295 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1296 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1297 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1298 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1299 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3544), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1300 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4700), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1301 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3544), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4700), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3670));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1302 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1303 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1304 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1305 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1306 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1307 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[45]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1308 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1310 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6900 (.Y(N12533), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6901 (.Y(N12523), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6902 (.Y(N12531), .A0(N12533), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652), .B0(N12523));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6903 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799), .A(N12531));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6826 (.Y(N12419), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6827 (.Y(N12420), .A(N12419));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1314 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806), .A(N12420));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1315 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[45]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[45]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1316 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1317 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1318 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3837), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1319 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3837));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1320 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4151), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1321 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3135), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1322 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3516), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3135), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1323 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4601), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3516));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1324 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4050), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1325 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3598), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1326 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4050), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3598));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1327 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[39]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4151), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4601), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1328 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1329 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3411), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1330 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[40]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3411));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1331 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1332 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[39]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[40]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1333 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1334 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1335 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4867), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1336 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3588), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1337 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3246), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3588));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1338 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[38]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4867), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3246), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1339 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[38]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[39]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1340 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1341 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1342 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3964), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1343 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3520), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1344 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[37]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3964), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3520), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1345 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[37]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[38]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1346 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4200), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1347 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[36]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4200), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1348 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[36]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[37]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1349 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1350 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7499), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1351 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1352 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1353 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4788), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1354 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4523), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1355 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3169), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4523));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1356 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[42]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4788), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3169), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1357 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1358 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1359 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4223), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1360 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3301), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1361 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3301));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1362 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4448), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4223), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1363 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4448));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1364 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1365 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1366 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[43]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819));
MXI2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1367 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[42]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[43]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1368 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[44]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[43]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1369 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7493), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[44]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1370 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1371 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1372 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4116), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1373 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4364), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1374 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4364));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1375 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4641), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4116), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1376 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4677), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4641));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1377 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4227), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1378 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[35]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4677), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4227), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1379 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[35]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[36]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1380 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1381 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1382 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4717), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1383 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3319), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4717));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1384 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4947), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1385 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[34]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3319), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4947), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1386 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[34]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[35]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1387 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1388 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1389 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3591), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1390 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4044), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1391 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[33]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3591), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4044), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6904 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803), .A0(N12533), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652), .B0(N12523));
INVXL buf1_A_I6934 (.Y(N12573), .A(N12531));
INVXL buf1_A_I6935 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47]), .A(N12573));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1393 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[33]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[34]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1394 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4997), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1395 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[32]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4997));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1396 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[32]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[33]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1397 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1398 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7532), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1399 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1400 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4825), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454));
INVXL buf1_A_I6828 (.Y(N12423), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915));
INVXL buf1_A_I6829 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006), .A(N12423));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1402 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4918), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718));
OAI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1403 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4375), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4918));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1404 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4825), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4375));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1405 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4355), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1406 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[30]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4355));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1407 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1408 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4306), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1409 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4753), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1410 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4306), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4753), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1411 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[30]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[31]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1412 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[31]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[32]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1413 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1414 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1415 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5025), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1416 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3402), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1417 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5103), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1418 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4651), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1419 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5103), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4651));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1420 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[29]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5025), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3402), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1421 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[29]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[30]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1422 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3721), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1423 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[28]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3721));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1424 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[28]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[29]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1425 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1426 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7433), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1427 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428), .A(N11299), .B(N11399));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1428 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1429 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3886), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1430 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3438), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1431 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[41]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3886), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3438), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1432 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[41]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[42]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1433 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[40]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[41]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1434 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41]));
NAND4BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1435 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7505), .AN(N11297), .B(N11368), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428), .D(N11372));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1436 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1437 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3672), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1438 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4118), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1439 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1440 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[27]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3672), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4118), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1441 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1442 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[27]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[28]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1443 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3080), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1444 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[26]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3080));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1445 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[26]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[27]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1446 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1447 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1448 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4831), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1449 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4384), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1450 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11836), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1451 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11836));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1452 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[25]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4831), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4384), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1453 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[25]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[26]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1454 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4512), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1455 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4512));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1456 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[24]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[25]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1457 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1458 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7467), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1459 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1460 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5096), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1461 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3482), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1462 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4091), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1463 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3434), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4091), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1464 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3434), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1465 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[23]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5096), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3482), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1466 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[23]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[24]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1467 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1468 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482), .A(N11401), .B(N10986));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1469 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1470 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7429), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7505), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1471 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3871), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1472 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3871), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1473 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22612), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[22]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[23]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1474 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663), .A(rm[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1475 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679), .A(rm[0]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1476 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22613), .A(rm[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1477 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788), .A(a_sign), .B(b_sign));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1478 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666), .A(rm[2]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1479 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684), .A(rm[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1480 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684));
AND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1481 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5), .A(rm[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1482 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1483 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22637), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22613), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1484 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22622), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1485 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1486 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3821), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1487 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4269), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1488 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1489 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3821), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4269), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1490 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1491 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1492 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3455), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1493 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3556), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3455));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1494 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3105), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1495 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3556), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3105), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1496 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802), .A(N12420));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1497 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[17]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[18]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1498 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4029), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1499 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4029));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1500 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[16]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[17]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1501 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7731), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[18]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[17]));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1502 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22569), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1503 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22579), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1504 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22563), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22579));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1505 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22569), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22563));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1506 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22560), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1507 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22560));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1508 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[14]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[15]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47]));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1509 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801), .A(N12420));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1510 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[15]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[16]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1511 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7742), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[15]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[16]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1512 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7751), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7742), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7731));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1513 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3479), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1514 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3479));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1515 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[13]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[14]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1516 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4187), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1517 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4187));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1518 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[12]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[13]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1519 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7753), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[14]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[13]));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1520 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4874), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1521 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4857), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4874), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1522 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4906), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1523 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4857), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4906));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1524 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[11]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[12]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1525 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3551), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1526 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3551));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1527 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[10]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[11]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1528 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7763), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[12]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[11]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1529 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7761), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7753), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7763));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1530 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22628), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7761));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1531 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1532 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5136), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1533 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5136));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1534 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[2]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1535 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807), .A(N12420));
OR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1536 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1537 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[0]), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[0]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1538 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[1]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1539 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7749), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[1]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1540 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7729), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7749));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1541 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1542 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3745), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1543 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4192), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1544 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3745), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4192), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1545 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[21]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[22]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1546 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3233), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1547 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3233));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1548 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[20]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[21]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1549 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7759), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[22]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[21]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1550 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1551 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1552 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5093), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1553 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3618), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1554 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3618));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1555 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3373), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5093), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1556 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4911), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1557 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4460), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1558 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4460), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1559 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[19]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[20]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1560 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[18]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[19]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1561 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7721), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[20]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[19]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1562 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7740), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7759), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7721));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1563 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7744), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7729), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7740));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1564 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3385), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1565 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4264), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865));
CLKXOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1566 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3385), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4264));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1567 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800), .A(N12420));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1568 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[10]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1569 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4985), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1570 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4985));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1571 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[9]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1572 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7725), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[10]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[9]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1573 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3630), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1574 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3630));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1575 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[8]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1576 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4341), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1577 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4341));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1578 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[7]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1579 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7735), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[7]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1580 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7723), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7725), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7735));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1581 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4423), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1582 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4423));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1583 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[3]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1584 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3708), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1585 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3708));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1586 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[4]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1587 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7757), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[4]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1588 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5062), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1589 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5062));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1590 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[6]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1591 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[5]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1592 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7746), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[5]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1593 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7733), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7757), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7746));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1594 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7738), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7723), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7733));
NAND3X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6933 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646), .A(N12110), .B(N12112), .C(N12147));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1597 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22619), .A(N10988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1598 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22615), .A(N11684), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22619));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1599 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22614), .A(N11658), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22615));
CLKBUFX3 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1600 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22617), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1601 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22631), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1602 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22641), .A(N11665), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22617));
OAI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1603 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44), .A0(N11646), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22614), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22641));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1604 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8524), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1605 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8524));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1606 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11903), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7429), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1607 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8421), .A(N10981), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11903));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1608 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3008), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1609 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3012), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1610 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3008), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3012));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1611 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2885), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1612 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2889), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1613 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2885), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2889));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1614 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13));
AND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1615 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__7), .A(rm[0]), .B(rm[1]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1616 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8254), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__7), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1617 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8254), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1618 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2919), .A(a_exp[7]), .B(a_exp[6]));
AND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1619 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2917), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1620 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11829), .A(a_exp[0]), .B(a_exp[1]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2917));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1621 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2919), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11829));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1622 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2955), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1623 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2959), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934), .B(a_man[0]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2955), .D(a_man[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1624 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2940), .A(a_man[10]), .B(a_man[9]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1625 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2961), .A(a_man[6]), .B(a_man[5]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1626 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2950), .A(a_man[8]), .B(a_man[7]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1627 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2971), .A(a_man[4]), .B(a_man[3]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1628 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2953), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2940), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2961), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2950), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2971));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1629 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2965), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1630 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2975), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1631 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2959), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2953), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2965), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2975));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1632 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1633 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2796), .A(b_exp[7]), .B(b_exp[6]));
AND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1634 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2794), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1635 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11821), .A(b_exp[0]), .B(b_exp[1]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2794));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1636 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2796), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11821));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1637 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2832), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1638 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2836), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811), .B(b_man[0]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2832), .D(b_man[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1639 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2817), .A(b_man[10]), .B(b_man[9]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1640 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2838), .A(b_man[6]), .B(b_man[5]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1641 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2827), .A(b_man[8]), .B(b_man[7]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1642 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2848), .A(b_man[4]), .B(b_man[3]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1643 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2830), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2817), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2838), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2827), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2848));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1644 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2842), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1645 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2852), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1646 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2836), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2830), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2842), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2852));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1647 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1648 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1649 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12));
AOI211XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1650 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3051), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22), .C0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1651 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3051));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1652 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1653 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8319), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1654 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857), .A(a_exp[7]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1655 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888), .A(b_exp[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1656 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7890), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1657 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852), .A(a_exp[6]), .B(b_exp[6]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1658 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897), .A(a_exp[5]), .B(b_exp[5]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1659 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1660 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861), .A(a_exp[4]), .B(b_exp[4]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1661 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908), .A(a_exp[3]), .B(b_exp[3]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1662 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1663 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7865), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1664 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870), .A(a_exp[2]), .B(b_exp[2]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1665 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916), .A(a_exp[1]), .B(b_exp[1]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1666 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7903), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1667 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879), .A(b_exp[0]), .B(a_exp[0]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1668 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900), .A(a_exp[1]), .B(b_exp[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1669 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854), .A(a_exp[2]), .B(b_exp[2]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1670 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7885), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1671 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7903), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7885));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1672 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892), .A(a_exp[3]), .B(b_exp[3]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1673 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920), .A(a_exp[4]), .B(b_exp[4]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1674 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1675 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881), .A(a_exp[5]), .B(b_exp[5]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1676 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913), .A(a_exp[6]), .B(b_exp[6]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1677 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7863), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1678 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7849), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7863));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1679 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7865), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7849));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1680 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867), .A(b_exp[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1681 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7869), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1682 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9]), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7890), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7869));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1683 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7915), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1684 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7899), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1685 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7915), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7899), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1686 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7868), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1687 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7868));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1688 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8228), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7]));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1689 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8228));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1690 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8319), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1691 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8507), .A(b_man[21]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1692 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8511), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8507), .B(a_man[21]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1693 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8545), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1694 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8545));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1695 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8467), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8511), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1696 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[8]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1697 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1698 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7864), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1699 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7923), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1700 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7907), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1701 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7891), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1702 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7907), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7891));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1703 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7864), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7923), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1704 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[6]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1705 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8015), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1706 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1707 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7918), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1708 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7904), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1709 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7918), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7904), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1710 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7878), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1711 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7878));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1712 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684), .A(b_exp[0]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1713 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696), .A(a_exp[0]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1714 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1715 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1716 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1717 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7902), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1718 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7902));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1719 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3]));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1720 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1721 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1722 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1723 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1724 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7874), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1725 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7895), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1726 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7874), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7895), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1727 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11840), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[4]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1728 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11840));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1729 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8015), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1730 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1731 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3390), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1732 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3095), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3390));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1733 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4711), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1734 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[46]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3095), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4711), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1735 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[47]), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[46]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1736 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[46]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[45]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[46]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1737 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1738 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22815), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1739 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22788), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22815), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1740 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22804), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1741 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22792), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22804), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1742 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22788), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22792));
AND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1743 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7506), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[47]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[46]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1744 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1745 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1746 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7540), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1747 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7534), .A(N12074), .B(N11377));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1748 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1749 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1750 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7473), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1751 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7469), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1752 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7486), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36]));
CLKAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1753 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441), .A(N12086), .B(N12091));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1754 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468), .A(N11462), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1755 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1756 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1757 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7511), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1758 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26]));
AND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1759 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1760 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1761 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495), .A(N12063), .B(N11464));
NOR3X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1762 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7534), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468));
AOI21X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6927 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[24]), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44), .B0(N11635));
CLKINVX6 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6928 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1765 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[8]), .A(N11528), .B(N11530), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1766 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1767 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[6]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1768 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8018), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1769 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8018), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1770 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[7]), .A(N11586), .B(N11584), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1771 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004));
MXI2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1772 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6]), .A(N11595), .B(N11593), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1773 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8136), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1774 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22677), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696), .B(a_exp[0]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1775 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681), .B(N11580));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1776 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6929 (.Y(N12555), .A(N11563));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6930 (.Y(N12551), .A(N11565));
MXI2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6931 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1]), .A(N12555), .B(N12551), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1778 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8132), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1]));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1779 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8130), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8136), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8132));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1780 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[4]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1781 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22861), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1782 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22856), .A(N11536), .B(N11538), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1783 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1784 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22871), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1785 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22869), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1786 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1787 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22865), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22869), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1788 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22872), .A(N11609), .B(N11607), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1789 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8140), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22856), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22872));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1790 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1791 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054), .A(N11554), .B(N11556), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1792 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8047), .A(N12025));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1793 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1794 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8047), .B(N11547), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1795 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8127), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3]));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1796 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8134), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8140), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8127));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1797 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8138), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8130), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8134));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1798 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7990), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1799 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8016), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1800 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8016));
MXI2XL mx2a_A_I6832 (.Y(N12434), .A(N11572), .B(N11574), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
INVXL mx2a_A_I6833 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9]), .A(N12434));
BUFX2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1802 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8157), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9]));
AOI21X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1803 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22706), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[8]), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8138), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8157));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1804 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[4]), .A(N11536), .B(N11538), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1805 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8176), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[8]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1806 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22987), .A(N11614), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1807 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[5]), .A(N11515), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22987));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1808 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[7]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1809 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8181), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1810 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8187), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8176), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8181));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1811 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8178), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[0]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1812 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8188), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1813 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8173), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1814 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8190), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8188), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8173));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1815 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8183), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8178), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8190));
OR3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1816 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8206), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1817 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8212), .A(N11360), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9]));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1818 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22693), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8187), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8183), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8212));
NOR2X4 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1819 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22685), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22706), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22693));
INVX12 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1820 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22685));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1821 (.Y(x[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8421), .B(N10691), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1822 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436), .A(N12063));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1823 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503), .A(N11462), .B(N11464));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1824 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7484), .A(N11377), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1825 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7551), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7484));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1826 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11896), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7551), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1827 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8374), .A(N10976), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11896));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1828 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8411), .A(b_man[20]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1829 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8463), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8411), .B(a_man[20]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1830 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8420), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8463), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1831 (.Y(x[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8374), .B(N10698), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1832 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7479), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1833 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7517), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1834 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7530), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1835 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470), .A(N12102));
CLKAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6834 (.Y(N12440), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6895 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6896 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550), .A(N12440));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I6897 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550));
NAND4BBXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1839 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7462), .AN(N11288), .BN(N11290), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470), .D(N12031));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1840 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[19]), .A(N11072), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7462));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1841 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8547), .A(N11072), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[19]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1842 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8536), .A(b_man[19]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1843 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8415), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8536), .B(a_man[19]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1844 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8371), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8415), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1845 (.Y(x[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8547), .B(N10705), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1846 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1847 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1848 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7520), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1849 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425), .A(N12084), .B(N12086));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1850 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1851 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7481), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1852 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455), .A(N12091), .B(N12096));
NAND4BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1853 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7512), .AN(N12123), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425), .C(N11143), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1854 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7512), .B(N11065));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1855 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8497), .A(N11065), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[18]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1856 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8442), .A(b_man[18]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1857 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8368), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8442), .B(a_man[18]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1858 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8543), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8368), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1859 (.Y(x[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8497), .B(N10712), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1860 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[0]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1861 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461), .A(N11399), .B(N11401));
NAND4BBXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1862 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7422), .AN(N11297), .BN(N11299), .C(N11293), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1863 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[17]), .A(N11058), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7422));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1864 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8452), .A(N11058), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[17]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1865 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8342), .A(b_man[17]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1866 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8539), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8342), .B(a_man[17]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1867 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8494), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8539), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1868 (.Y(x[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8452), .B(N10719), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1869 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7439), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1870 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11889), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7439), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1871 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8403), .A(N10971), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11889));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1872 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8468), .A(b_man[16]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1873 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8489), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8468), .B(a_man[16]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1874 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8450), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8489), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1875 (.Y(x[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8403), .B(N10726), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1876 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7543), .A(N12081), .B(N12418));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1877 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524), .A(N12100), .B(N12102));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1878 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7459), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7543), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1879 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7459), .B(N11051));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1880 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8352), .A(N11051), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[15]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1881 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8373), .A(b_man[15]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1882 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8373), .B(a_man[15]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1883 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8400), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8446), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1884 (.Y(x[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8352), .B(N10733), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1885 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455), .B(N11418));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1886 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7437), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1887 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7432), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485), .B(N12119));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1888 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7432), .B(N11044));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1889 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8526), .A(N11044), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[14]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1890 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8495), .A(b_man[14]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1891 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8396), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8495), .B(a_man[14]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1892 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8351), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8396), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1893 (.Y(x[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8526), .B(N10740), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1894 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7537), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1895 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7537), .B(N11037));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1896 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8477), .A(N11037), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[13]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1897 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8401), .A(b_man[13]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1898 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8346), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8401), .B(a_man[13]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1899 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8522), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8346), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1900 (.Y(x[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8477), .B(N10747), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1901 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7508), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503), .B(N12063));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1902 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7508), .B(N11030));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1903 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8432), .A(N11030), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[12]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1904 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8525), .A(b_man[12]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1905 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8519), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8525), .B(a_man[12]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1906 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8474), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8519), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1907 (.Y(x[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8432), .B(N10754), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1908 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7476), .A(N12031), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1909 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7476), .B(N11023));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1910 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8383), .A(N11023), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[11]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1911 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8430), .A(b_man[11]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1912 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8470), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8430), .B(a_man[11]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1913 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8429), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8470), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1914 (.Y(x[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8383), .B(N10761), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1915 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7491), .A(N12123), .B(N11304));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1916 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11882), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7491), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1917 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8556), .A(N10966), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11882));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1918 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8554), .A(b_man[10]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1919 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8423), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8554), .B(a_man[10]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1920 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8381), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8423), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1921 (.Y(x[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8556), .B(N10768), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1922 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7475), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461), .B(N11293));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1923 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7475), .B(N11016));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1924 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8506), .A(N11016), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[9]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1925 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8458), .A(b_man[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1926 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8377), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8458), .B(a_man[9]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1927 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8553), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8377), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1928 (.Y(x[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8506), .B(N10775), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1929 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495), .B(N11009));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1930 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8459), .A(N11009), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[8]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1931 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8361), .A(b_man[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1932 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8549), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8361), .B(a_man[8]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1933 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8504), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8549), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1934 (.Y(x[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8459), .B(N10782), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1935 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11875), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1936 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8410), .A(N10961), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11875));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1937 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8484), .A(b_man[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1938 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8499), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8484), .B(a_man[7]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1939 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8457), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8499), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1940 (.Y(x[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8410), .B(N10789), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1941 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494), .A(N12119));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1942 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11868), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1943 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8363), .A(N10956), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11868));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1944 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8390), .A(b_man[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1945 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8454), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8390), .B(a_man[6]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1946 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8408), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8454), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1947 (.Y(x[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8363), .B(N10796), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1948 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464), .B(N11002));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1949 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8535), .A(N11002), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[5]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1950 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8512), .A(b_man[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1951 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8404), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8512), .B(a_man[5]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1952 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8360), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8404), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1953 (.Y(x[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8535), .B(N10803), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1954 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436), .B(N10995));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1955 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8486), .A(N10995), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[4]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1956 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8417), .A(b_man[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1957 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8354), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8417), .B(a_man[4]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1958 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8533), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8354), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1959 (.Y(x[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8486), .B(N10810), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1960 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11861), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1961 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8440), .A(N10951), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11861));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1962 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8541), .A(b_man[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1963 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8529), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8541), .B(a_man[3]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1964 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8483), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8529), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1965 (.Y(x[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8440), .B(N10817), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1966 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11854), .A(N11143), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1967 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8391), .A(N10946), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11854));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1968 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8447), .A(b_man[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1969 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8479), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8447), .B(a_man[2]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1970 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8439), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8479), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1971 (.Y(x[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8391), .B(N10824), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1972 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11847), .A(N11293), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1973 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8341), .A(N10941), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11847));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1974 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8348), .A(b_man[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1975 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8434), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8348), .B(a_man[1]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1976 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8388), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8434), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1977 (.Y(x[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8341), .B(N10831), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1978 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8515), .A(N10988), .B(N10986), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1979 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8472), .A(b_man[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1980 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8384), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8472), .B(a_man[0]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1981 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8337), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8384), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1982 (.Y(x[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8515), .B(N10838), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1983 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7522), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435));
NAND4BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1984 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7456), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485), .B(N11261), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1985 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7456), .B(N11079));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1986 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8324), .A(N11079), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[22]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1987 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8329), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1988 (.Y(x[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8324), .B(N12104), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1989 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1990 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8288), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1991 (.Y(x[30]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861), .B(N10852), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1992 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8282), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1993 (.Y(x[29]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8282), .B(N10852), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1994 (.Y(x[28]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[5]), .B(N10852), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1995 (.Y(x[27]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[4]), .B(N10852), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1996 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8263), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1997 (.Y(x[26]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8263), .B(N10852), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1998 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8285), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I1999 (.Y(x[25]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8285), .B(N10852), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2000 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8279), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2001 (.Y(x[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8279), .B(N10852), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2002 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22682), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38), .S0(N11100));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2003 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22689), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469));
NOR3XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2004 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22678), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22689), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2005 (.Y(x[23]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22682), .B(N10901), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2006 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3068), .AN(b_sign), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2007 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3074), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3068), .B(a_sign), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_2_I2008 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3074), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26));
reg x_reg_31__I2040_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I2040_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[31];
	end
assign x[31] = x_reg_31__I2040_QOUT;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[44] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[23] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[0] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[4] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[5] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[1] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[2] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[3] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[6] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[7] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[10] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[16] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[20] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[21] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[23] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[2] = 1'B0;
endmodule

/* CADENCE  s7P5SA3eqhw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



