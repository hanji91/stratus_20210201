/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:28 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_5 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456;
wire N4120,N8900,N8938,N8945,N8952,N8958,N8961 
	,N8970,N8979,N8988,N8997,N9006,N9015,N9024,N9033 
	,N9042,N9051,N9060,N9069,N9078,N9087,N9096,N9105 
	,N9114,N9123,N9132,N9141,N9152,N9157,N9162,N9167 
	,N9172,N9177,N9182,N9187,N9192,N9197,N9202,N9207 
	,N9212,N9217,N9222,N9227,N9232,N9237,N9242,N9247 
	,N9252,N9257,N9624,N9631,N9633,N9638,N9645,N9652 
	,N9659,N9666,N9671,N9673,N9678,N9680,N9706,N9732 
	,N9758,N9925,N9931,N9934,N9943,N9952,N9961,N9970 
	,N9979,N9988,N9997,N10006,N10015,N10024,N10033,N10042 
	,N10051,N10060,N10069,N10078,N10087,N10096,N10105,N10114 
	,N10125,N10130,N10135,N10140,N10145,N10150,N10155,N10160 
	,N10165,N10170,N10175,N10180,N10185,N10190,N10195,N10200 
	,N10205,N10210,N10215,N10220,N10225,N10230,N10233,N10239 
	,N10242,N10248,N10251,N10257,N10260,N10266,N10269,N10275 
	,N10278,N10284,N10287,N10293,N10296,N10302,N10305,N10311 
	,N10314,N10320,N10323,N10329,N10332,N10338,N10341,N10347 
	,N10350,N10356,N10359,N10365,N10368,N10374,N10377,N10383 
	,N10386,N10392,N10395,N10401,N10404,N10410,N10413,N10419 
	,N10422,N10428,N10567,N10593,N10619,N10645,N10751,N10753 
	,N10790,N10792,N10798,N10800,N10812,N10814,N10821,N10823 
	,N10830,N10832,N10839,N10841,N10858,N10860,N10867,N10869 
	,N10876,N10878,N10885,N10887,N10921,N10923,N10925,N10969 
	,N10971,N10973,N11301,N11307,N11313,N11319,N11325,N11331 
	,N11337,N11343,N11349,N11355,N11361,N11451,N11453,N11458 
	,N11460,N11465,N11467,N11472,N11479,N11481,N11488,N11495 
	,N11500,N11502,N11507,N11521,N11523,N11536,N11539,N11549 
	,N11552,N11559,N11566,N11573,N11583,N11589,N11592,N11610 
	,N11624,N11643,N11645,N11658,N11662,N11664,N11672,N11678 
	,N11684,N11692,N11694,N11702,N11710,N11712,N11717,N11727 
	,N11733,N11739,N11742,N11752,N11756,N11758,N11791,N11793 
	,N11802,N11804,N11810,N11812,N11821,N11823,N11829,N11831 
	,N11835,N11837,N11840,N11904,N11906,N11930,N11941,N11949 
	,N11951,N11960,N11962,N11971,N11973,N11981,N11983,N12644 
	,N12649,N12652,N12655,N12658,N12662,N13247,N13248,N13249 
	,N13250,N13251,N13252,N13253,N13254,N13255,N13256,N13257 
	,N13258,N13259,N13260,N13261,N13262,N13263,N13264,N13265 
	,N13266,N13267,N13268,N13270,N13271,N13273,N13280,N13287 
	,N13294,N13303,N13309,N13311,N13319;
reg x_reg_L1_21__retimed_I6582_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I6582_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49;
	end
assign N12662 = x_reg_L1_21__retimed_I6582_QOUT;
assign N13247 = !N12662;
assign N13248 = !N13247;
reg x_reg_L0_21__retimed_I6580_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6580_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384;
	end
assign N12658 = x_reg_L0_21__retimed_I6580_QOUT;
reg x_reg_L0_21__retimed_I6579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6579_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751;
	end
assign N12655 = x_reg_L0_21__retimed_I6579_QOUT;
reg x_reg_L0_21__retimed_I6578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6578_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275;
	end
assign N12652 = x_reg_L0_21__retimed_I6578_QOUT;
reg x_reg_L0_21__retimed_I6577_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6577_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613;
	end
assign N12649 = x_reg_L0_21__retimed_I6577_QOUT;
reg x_reg_L0_21__retimed_I6575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6575_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[20];
	end
assign N12644 = x_reg_L0_21__retimed_I6575_QOUT;
reg x_reg_L0_21__retimed_I6291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6291_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922;
	end
assign N11983 = x_reg_L0_21__retimed_I6291_QOUT;
reg x_reg_L0_21__retimed_I6290_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6290_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563;
	end
assign N11981 = x_reg_L0_21__retimed_I6290_QOUT;
reg x_reg_L0_21__retimed_I6288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6288_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016;
	end
assign N11973 = x_reg_L0_21__retimed_I6288_QOUT;
reg x_reg_L0_21__retimed_I6287_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6287_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651;
	end
assign N11971 = x_reg_L0_21__retimed_I6287_QOUT;
reg x_reg_L0_21__retimed_I6284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6284_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501;
	end
assign N11962 = x_reg_L0_21__retimed_I6284_QOUT;
reg x_reg_L0_21__retimed_I6283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6283_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099;
	end
assign N11960 = x_reg_L0_21__retimed_I6283_QOUT;
reg x_reg_L0_21__retimed_I6280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6280_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415;
	end
assign N11951 = x_reg_L0_21__retimed_I6280_QOUT;
reg x_reg_L0_21__retimed_I6279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6279_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342;
	end
assign N11949 = x_reg_L0_21__retimed_I6279_QOUT;
reg x_reg_L0_21__retimed_I6276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6276_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811;
	end
assign N11941 = x_reg_L0_21__retimed_I6276_QOUT;
reg x_reg_L0_21__retimed_I6272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6272_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244;
	end
assign N11930 = x_reg_L0_21__retimed_I6272_QOUT;
reg x_reg_L0_21__retimed_I6264_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6264_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824;
	end
assign N11906 = x_reg_L0_21__retimed_I6264_QOUT;
reg x_reg_L0_21__retimed_I6263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6263_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185;
	end
assign N11904 = x_reg_L0_21__retimed_I6263_QOUT;
reg x_reg_L0_21__retimed_I6257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6257_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656;
	end
assign N11840 = x_reg_L0_21__retimed_I6257_QOUT;
reg x_reg_L0_21__retimed_I6256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6256_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314;
	end
assign N11837 = x_reg_L0_21__retimed_I6256_QOUT;
reg x_reg_L0_21__retimed_I6255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6255_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495;
	end
assign N11835 = x_reg_L0_21__retimed_I6255_QOUT;
reg x_reg_L0_21__retimed_I6254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6254_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396;
	end
assign N11831 = x_reg_L0_21__retimed_I6254_QOUT;
reg x_reg_L0_21__retimed_I6253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6253_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471;
	end
assign N11829 = x_reg_L0_21__retimed_I6253_QOUT;
reg x_reg_L0_21__retimed_I6251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6251_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694;
	end
assign N11823 = x_reg_L0_21__retimed_I6251_QOUT;
reg x_reg_L0_21__retimed_I6250_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6250_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435;
	end
assign N11821 = x_reg_L0_21__retimed_I6250_QOUT;
reg x_reg_L0_21__retimed_I6247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6247_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413;
	end
assign N11812 = x_reg_L0_21__retimed_I6247_QOUT;
reg x_reg_L0_21__retimed_I6246_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6246_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073;
	end
assign N11810 = x_reg_L0_21__retimed_I6246_QOUT;
reg x_reg_L0_21__retimed_I6244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6244_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171;
	end
assign N11804 = x_reg_L0_21__retimed_I6244_QOUT;
reg x_reg_L0_21__retimed_I6243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6243_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524;
	end
assign N11802 = x_reg_L0_21__retimed_I6243_QOUT;
reg x_reg_L0_21__retimed_I6240_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6240_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669;
	end
assign N11793 = x_reg_L0_21__retimed_I6240_QOUT;
reg x_reg_L0_21__retimed_I6239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6239_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036;
	end
assign N11791 = x_reg_L0_21__retimed_I6239_QOUT;
reg x_reg_L0_21__retimed_I6225_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6225_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539;
	end
assign N11758 = x_reg_L0_21__retimed_I6225_QOUT;
reg x_reg_L0_21__retimed_I6224_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6224_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185;
	end
assign N11756 = x_reg_L0_21__retimed_I6224_QOUT;
reg x_reg_L0_21__retimed_I6223_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6223_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112;
	end
assign N11752 = x_reg_L0_21__retimed_I6223_QOUT;
reg x_reg_L0_21__retimed_I6219_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6219_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256;
	end
assign N11742 = x_reg_L0_21__retimed_I6219_QOUT;
reg x_reg_L0_21__retimed_I6218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6218_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193;
	end
assign N11739 = x_reg_L0_21__retimed_I6218_QOUT;
reg x_reg_L0_21__retimed_I6216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6216_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904;
	end
assign N11733 = x_reg_L0_21__retimed_I6216_QOUT;
reg x_reg_L0_21__retimed_I6214_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6214_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596;
	end
assign N11727 = x_reg_L0_21__retimed_I6214_QOUT;
reg x_reg_L0_21__retimed_I6210_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6210_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423;
	end
assign N11717 = x_reg_L0_21__retimed_I6210_QOUT;
reg x_reg_L0_21__retimed_I6208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6208_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733;
	end
assign N11712 = x_reg_L0_21__retimed_I6208_QOUT;
reg x_reg_L0_21__retimed_I6207_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6207_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389;
	end
assign N11710 = x_reg_L0_21__retimed_I6207_QOUT;
reg x_reg_L0_21__retimed_I6205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6205_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197;
	end
assign N11702 = x_reg_L0_21__retimed_I6205_QOUT;
reg x_reg_L0_21__retimed_I6202_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6202_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527;
	end
assign N11694 = x_reg_L0_21__retimed_I6202_QOUT;
reg x_reg_L0_21__retimed_I6201_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6201_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191;
	end
assign N11692 = x_reg_L0_21__retimed_I6201_QOUT;
reg x_reg_L0_21__retimed_I6199_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6199_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787;
	end
assign N11684 = x_reg_L0_21__retimed_I6199_QOUT;
reg x_reg_L0_21__retimed_I6197_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6197_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274;
	end
assign N11678 = x_reg_L0_21__retimed_I6197_QOUT;
reg x_reg_L0_21__retimed_I6195_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6195_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995;
	end
assign N11672 = x_reg_L0_21__retimed_I6195_QOUT;
reg x_reg_L0_21__retimed_I6192_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6192_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333;
	end
assign N11664 = x_reg_L0_21__retimed_I6192_QOUT;
reg x_reg_L0_21__retimed_I6191_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6191_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986;
	end
assign N11662 = x_reg_L0_21__retimed_I6191_QOUT;
reg x_reg_L0_21__retimed_I6190_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6190_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680;
	end
assign N11658 = x_reg_L0_21__retimed_I6190_QOUT;
reg x_reg_L0_21__retimed_I6185_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6185_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[18];
	end
assign N11645 = x_reg_L0_21__retimed_I6185_QOUT;
reg x_reg_L0_21__retimed_I6184_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6184_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[17];
	end
assign N11643 = x_reg_L0_21__retimed_I6184_QOUT;
reg x_reg_L0_21__retimed_I6176_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6176_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[19];
	end
assign N11624 = x_reg_L0_21__retimed_I6176_QOUT;
reg x_reg_L0_21__retimed_I6170_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6170_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[0];
	end
assign N11610 = x_reg_L0_21__retimed_I6170_QOUT;
reg x_reg_L0_21__retimed_I6162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6162_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055;
	end
assign N11592 = x_reg_L0_21__retimed_I6162_QOUT;
reg x_reg_L0_21__retimed_I6161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6161_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395;
	end
assign N11589 = x_reg_L0_21__retimed_I6161_QOUT;
reg x_reg_L0_21__retimed_I6159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6159_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692;
	end
assign N11583 = x_reg_L0_21__retimed_I6159_QOUT;
reg x_reg_L0_21__retimed_I6155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6155_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219;
	end
assign N11573 = x_reg_L0_21__retimed_I6155_QOUT;
reg x_reg_L0_21__retimed_I6152_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6152_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623;
	end
assign N11566 = x_reg_L0_21__retimed_I6152_QOUT;
reg x_reg_L0_21__retimed_I6149_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6149_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422;
	end
assign N11559 = x_reg_L0_21__retimed_I6149_QOUT;
reg x_reg_L0_21__retimed_I6146_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6146_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225;
	end
assign N11552 = x_reg_L0_21__retimed_I6146_QOUT;
reg x_reg_L0_21__retimed_I6145_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6145_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571;
	end
assign N11549 = x_reg_L0_21__retimed_I6145_QOUT;
reg x_reg_L0_21__retimed_I6141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6141_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025;
	end
assign N11539 = x_reg_L0_21__retimed_I6141_QOUT;
reg x_reg_L0_21__retimed_I6140_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6140_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480;
	end
assign N11536 = x_reg_L0_21__retimed_I6140_QOUT;
reg x_reg_L0_21__retimed_I6135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6135_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[16];
	end
assign N11523 = x_reg_L0_21__retimed_I6135_QOUT;
reg x_reg_L0_21__retimed_I6134_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6134_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[15];
	end
assign N11521 = x_reg_L0_21__retimed_I6134_QOUT;
reg x_reg_L0_21__retimed_I6128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6128_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[3];
	end
assign N11507 = x_reg_L0_21__retimed_I6128_QOUT;
reg x_reg_L0_21__retimed_I6126_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6126_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[12];
	end
assign N11502 = x_reg_L0_21__retimed_I6126_QOUT;
reg x_reg_L0_21__retimed_I6125_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6125_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[11];
	end
assign N11500 = x_reg_L0_21__retimed_I6125_QOUT;
reg x_reg_L0_21__retimed_I6123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6123_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[7];
	end
assign N11495 = x_reg_L0_21__retimed_I6123_QOUT;
reg x_reg_L0_21__retimed_I6120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6120_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[6];
	end
assign N11488 = x_reg_L0_21__retimed_I6120_QOUT;
reg x_reg_L0_21__retimed_I6117_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6117_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[14];
	end
assign N11481 = x_reg_L0_21__retimed_I6117_QOUT;
reg x_reg_L0_21__retimed_I6116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6116_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[13];
	end
assign N11479 = x_reg_L0_21__retimed_I6116_QOUT;
reg x_reg_L0_21__retimed_I6113_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6113_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[8];
	end
assign N11472 = x_reg_L0_21__retimed_I6113_QOUT;
reg x_reg_L0_21__retimed_I6111_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6111_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[2];
	end
assign N11467 = x_reg_L0_21__retimed_I6111_QOUT;
reg x_reg_L0_21__retimed_I6110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6110_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[1];
	end
assign N11465 = x_reg_L0_21__retimed_I6110_QOUT;
reg x_reg_L0_21__retimed_I6108_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6108_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[10];
	end
assign N11460 = x_reg_L0_21__retimed_I6108_QOUT;
reg x_reg_L0_21__retimed_I6107_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6107_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[9];
	end
assign N11458 = x_reg_L0_21__retimed_I6107_QOUT;
reg x_reg_L0_21__retimed_I6105_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6105_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[5];
	end
assign N11453 = x_reg_L0_21__retimed_I6105_QOUT;
reg x_reg_L0_21__retimed_I6104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6104_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[4];
	end
assign N11451 = x_reg_L0_21__retimed_I6104_QOUT;
reg x_reg_L0_21__retimed_I6073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6073_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483;
	end
assign N11361 = x_reg_L0_21__retimed_I6073_QOUT;
reg x_reg_L0_21__retimed_I6071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6071_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360;
	end
assign N11355 = x_reg_L0_21__retimed_I6071_QOUT;
reg x_reg_L0_21__retimed_I6069_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6069_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161;
	end
assign N11349 = x_reg_L0_21__retimed_I6069_QOUT;
reg x_reg_L0_21__retimed_I6067_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6067_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564;
	end
assign N11343 = x_reg_L0_21__retimed_I6067_QOUT;
reg x_reg_L0_21__retimed_I6065_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6065_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284;
	end
assign N11337 = x_reg_L0_21__retimed_I6065_QOUT;
reg x_reg_L0_21__retimed_I6063_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6063_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082;
	end
assign N11331 = x_reg_L0_21__retimed_I6063_QOUT;
reg x_reg_L0_21__retimed_I6061_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6061_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367;
	end
assign N11325 = x_reg_L0_21__retimed_I6061_QOUT;
reg x_reg_L0_21__retimed_I6059_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6059_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166;
	end
assign N11319 = x_reg_L0_21__retimed_I6059_QOUT;
reg x_reg_L0_21__retimed_I6057_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6057_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869;
	end
assign N11313 = x_reg_L0_21__retimed_I6057_QOUT;
reg x_reg_L0_21__retimed_I6055_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6055_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659;
	end
assign N11307 = x_reg_L0_21__retimed_I6055_QOUT;
reg x_reg_L0_21__retimed_I6053_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6053_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449;
	end
assign N11301 = x_reg_L0_21__retimed_I6053_QOUT;
reg x_reg_L0_21__retimed_I5946_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5946_QOUT <= rm[2];
	end
assign N10973 = x_reg_L0_21__retimed_I5946_QOUT;
reg x_reg_L0_21__retimed_I5945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5945_QOUT <= rm[0];
	end
assign N10971 = x_reg_L0_21__retimed_I5945_QOUT;
reg x_reg_L0_21__retimed_I5944_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5944_QOUT <= rm[1];
	end
assign N10969 = x_reg_L0_21__retimed_I5944_QOUT;
reg x_reg_L0_21__retimed_I5929_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5929_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446;
	end
assign N10925 = x_reg_L0_21__retimed_I5929_QOUT;
reg x_reg_L0_21__retimed_I5928_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5928_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445;
	end
assign N10923 = x_reg_L0_21__retimed_I5928_QOUT;
reg x_reg_L0_21__retimed_I5927_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5927_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N10921 = x_reg_L0_21__retimed_I5927_QOUT;
reg x_reg_L0_21__retimed_I5918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5918_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3];
	end
assign N10887 = x_reg_L0_21__retimed_I5918_QOUT;
reg x_reg_L0_21__retimed_I5917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5917_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[3];
	end
assign N10885 = x_reg_L0_21__retimed_I5917_QOUT;
reg x_reg_L0_21__retimed_I5915_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5915_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7];
	end
assign N10878 = x_reg_L0_21__retimed_I5915_QOUT;
reg x_reg_L0_21__retimed_I5914_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5914_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[7];
	end
assign N10876 = x_reg_L0_21__retimed_I5914_QOUT;
reg x_reg_L0_21__retimed_I5912_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5912_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4];
	end
assign N10869 = x_reg_L0_21__retimed_I5912_QOUT;
reg x_reg_L0_21__retimed_I5911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5911_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[4];
	end
assign N10867 = x_reg_L0_21__retimed_I5911_QOUT;
reg x_reg_L0_21__retimed_I5909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5909_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2];
	end
assign N10860 = x_reg_L0_21__retimed_I5909_QOUT;
reg x_reg_L0_21__retimed_I5908_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5908_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[2];
	end
assign N10858 = x_reg_L0_21__retimed_I5908_QOUT;
reg x_reg_L0_21__retimed_I5902_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5902_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1];
	end
assign N10841 = x_reg_L0_21__retimed_I5902_QOUT;
reg x_reg_L0_21__retimed_I5901_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5901_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[1];
	end
assign N10839 = x_reg_L0_21__retimed_I5901_QOUT;
reg x_reg_L0_21__retimed_I5899_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5899_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6];
	end
assign N10832 = x_reg_L0_21__retimed_I5899_QOUT;
reg x_reg_L0_21__retimed_I5898_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5898_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[6];
	end
assign N10830 = x_reg_L0_21__retimed_I5898_QOUT;
reg x_reg_L0_21__retimed_I5896_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5896_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5];
	end
assign N10823 = x_reg_L0_21__retimed_I5896_QOUT;
reg x_reg_L0_21__retimed_I5895_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5895_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[5];
	end
assign N10821 = x_reg_L0_21__retimed_I5895_QOUT;
reg x_reg_L0_21__retimed_I5893_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5893_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0];
	end
assign N10814 = x_reg_L0_21__retimed_I5893_QOUT;
reg x_reg_L0_21__retimed_I5892_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5892_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0];
	end
assign N10812 = x_reg_L0_21__retimed_I5892_QOUT;
reg x_reg_L0_21__retimed_I5888_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5888_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8];
	end
assign N10800 = x_reg_L0_21__retimed_I5888_QOUT;
reg x_reg_L0_21__retimed_I5887_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5887_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[8];
	end
assign N10798 = x_reg_L0_21__retimed_I5887_QOUT;
reg x_reg_L0_21__retimed_I5885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5885_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9];
	end
assign N10792 = x_reg_L0_21__retimed_I5885_QOUT;
reg x_reg_L0_21__retimed_I5884_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5884_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[9];
	end
assign N10790 = x_reg_L0_21__retimed_I5884_QOUT;
reg x_reg_L0_21__retimed_I5869_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5869_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27;
	end
assign N10753 = x_reg_L0_21__retimed_I5869_QOUT;
reg x_reg_L0_21__retimed_I5868_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5868_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28;
	end
assign N10751 = x_reg_L0_21__retimed_I5868_QOUT;
reg x_reg_L1_21__retimed_I5842_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5842_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44;
	end
assign N10645 = x_reg_L1_21__retimed_I5842_QOUT;
reg x_reg_L1_21__retimed_I5840_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5840_QOUT <= N9758;
	end
assign N10619 = x_reg_L1_21__retimed_I5840_QOUT;
reg x_reg_L1_21__retimed_I5838_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5838_QOUT <= N9732;
	end
assign N10593 = x_reg_L1_21__retimed_I5838_QOUT;
reg x_reg_L1_21__retimed_I5836_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5836_QOUT <= N9706;
	end
assign N10567 = x_reg_L1_21__retimed_I5836_QOUT;
reg x_reg_L1_21__retimed_I5789_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5789_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45];
	end
assign N10428 = x_reg_L1_21__retimed_I5789_QOUT;
reg x_reg_L1_21__retimed_I5786_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5786_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[21];
	end
assign N10422 = x_reg_L1_21__retimed_I5786_QOUT;
reg x_reg_L1_20__retimed_I5785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5785_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44];
	end
assign N10419 = x_reg_L1_20__retimed_I5785_QOUT;
reg x_reg_L1_20__retimed_I5782_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5782_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[20];
	end
assign N10413 = x_reg_L1_20__retimed_I5782_QOUT;
reg x_reg_L1_19__retimed_I5781_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5781_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43];
	end
assign N10410 = x_reg_L1_19__retimed_I5781_QOUT;
reg x_reg_L1_19__retimed_I5778_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5778_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[19];
	end
assign N10404 = x_reg_L1_19__retimed_I5778_QOUT;
reg x_reg_L1_18__retimed_I5777_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5777_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42];
	end
assign N10401 = x_reg_L1_18__retimed_I5777_QOUT;
reg x_reg_L1_18__retimed_I5774_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5774_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[18];
	end
assign N10395 = x_reg_L1_18__retimed_I5774_QOUT;
reg x_reg_L1_17__retimed_I5773_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5773_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41];
	end
assign N10392 = x_reg_L1_17__retimed_I5773_QOUT;
reg x_reg_L1_17__retimed_I5770_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5770_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[17];
	end
assign N10386 = x_reg_L1_17__retimed_I5770_QOUT;
reg x_reg_L1_16__retimed_I5769_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5769_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40];
	end
assign N10383 = x_reg_L1_16__retimed_I5769_QOUT;
reg x_reg_L1_16__retimed_I5766_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5766_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[16];
	end
assign N10377 = x_reg_L1_16__retimed_I5766_QOUT;
reg x_reg_L1_15__retimed_I5765_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5765_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39];
	end
assign N10374 = x_reg_L1_15__retimed_I5765_QOUT;
reg x_reg_L1_15__retimed_I5762_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5762_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[15];
	end
assign N10368 = x_reg_L1_15__retimed_I5762_QOUT;
reg x_reg_L1_14__retimed_I5761_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5761_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38];
	end
assign N10365 = x_reg_L1_14__retimed_I5761_QOUT;
reg x_reg_L1_14__retimed_I5758_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5758_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[14];
	end
assign N10359 = x_reg_L1_14__retimed_I5758_QOUT;
reg x_reg_L1_13__retimed_I5757_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5757_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37];
	end
assign N10356 = x_reg_L1_13__retimed_I5757_QOUT;
reg x_reg_L1_13__retimed_I5754_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5754_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[13];
	end
assign N10350 = x_reg_L1_13__retimed_I5754_QOUT;
reg x_reg_L1_12__retimed_I5753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5753_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36];
	end
assign N10347 = x_reg_L1_12__retimed_I5753_QOUT;
reg x_reg_L1_12__retimed_I5750_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5750_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[12];
	end
assign N10341 = x_reg_L1_12__retimed_I5750_QOUT;
reg x_reg_L1_11__retimed_I5749_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5749_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35];
	end
assign N10338 = x_reg_L1_11__retimed_I5749_QOUT;
reg x_reg_L1_11__retimed_I5746_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5746_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[11];
	end
assign N10332 = x_reg_L1_11__retimed_I5746_QOUT;
reg x_reg_L1_10__retimed_I5745_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5745_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34];
	end
assign N10329 = x_reg_L1_10__retimed_I5745_QOUT;
reg x_reg_L1_10__retimed_I5742_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5742_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[10];
	end
assign N10323 = x_reg_L1_10__retimed_I5742_QOUT;
reg x_reg_L1_9__retimed_I5741_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5741_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33];
	end
assign N10320 = x_reg_L1_9__retimed_I5741_QOUT;
reg x_reg_L1_9__retimed_I5738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5738_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[9];
	end
assign N10314 = x_reg_L1_9__retimed_I5738_QOUT;
reg x_reg_L1_8__retimed_I5737_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5737_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32];
	end
assign N10311 = x_reg_L1_8__retimed_I5737_QOUT;
reg x_reg_L1_8__retimed_I5734_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5734_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[8];
	end
assign N10305 = x_reg_L1_8__retimed_I5734_QOUT;
reg x_reg_L1_7__retimed_I5733_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5733_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31];
	end
assign N10302 = x_reg_L1_7__retimed_I5733_QOUT;
reg x_reg_L1_7__retimed_I5730_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5730_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[7];
	end
assign N10296 = x_reg_L1_7__retimed_I5730_QOUT;
reg x_reg_L1_6__retimed_I5729_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5729_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30];
	end
assign N10293 = x_reg_L1_6__retimed_I5729_QOUT;
reg x_reg_L1_6__retimed_I5726_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5726_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[6];
	end
assign N10287 = x_reg_L1_6__retimed_I5726_QOUT;
reg x_reg_L1_5__retimed_I5725_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5725_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29];
	end
assign N10284 = x_reg_L1_5__retimed_I5725_QOUT;
reg x_reg_L1_5__retimed_I5722_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5722_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[5];
	end
assign N10278 = x_reg_L1_5__retimed_I5722_QOUT;
reg x_reg_L1_4__retimed_I5721_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5721_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28];
	end
assign N10275 = x_reg_L1_4__retimed_I5721_QOUT;
reg x_reg_L1_4__retimed_I5718_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5718_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[4];
	end
assign N10269 = x_reg_L1_4__retimed_I5718_QOUT;
reg x_reg_L1_3__retimed_I5717_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5717_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27];
	end
assign N10266 = x_reg_L1_3__retimed_I5717_QOUT;
reg x_reg_L1_3__retimed_I5714_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5714_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[3];
	end
assign N10260 = x_reg_L1_3__retimed_I5714_QOUT;
reg x_reg_L1_2__retimed_I5713_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5713_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26];
	end
assign N10257 = x_reg_L1_2__retimed_I5713_QOUT;
reg x_reg_L1_2__retimed_I5710_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5710_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N10251 = x_reg_L1_2__retimed_I5710_QOUT;
reg x_reg_L1_1__retimed_I5709_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5709_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25];
	end
assign N10248 = x_reg_L1_1__retimed_I5709_QOUT;
reg x_reg_L1_1__retimed_I5706_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5706_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N10242 = x_reg_L1_1__retimed_I5706_QOUT;
reg x_reg_L1_0__retimed_I5705_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5705_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24];
	end
assign N10239 = x_reg_L1_0__retimed_I5705_QOUT;
reg x_reg_L1_0__retimed_I5702_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5702_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N10233 = x_reg_L1_0__retimed_I5702_QOUT;
reg x_reg_L1_21__retimed_I5701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5701_QOUT <= N9257;
	end
assign N10230 = x_reg_L1_21__retimed_I5701_QOUT;
reg x_reg_L1_20__retimed_I5699_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5699_QOUT <= N9252;
	end
assign N10225 = x_reg_L1_20__retimed_I5699_QOUT;
reg x_reg_L1_19__retimed_I5697_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5697_QOUT <= N9247;
	end
assign N10220 = x_reg_L1_19__retimed_I5697_QOUT;
reg x_reg_L1_18__retimed_I5695_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5695_QOUT <= N9242;
	end
assign N10215 = x_reg_L1_18__retimed_I5695_QOUT;
reg x_reg_L1_17__retimed_I5693_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5693_QOUT <= N9237;
	end
assign N10210 = x_reg_L1_17__retimed_I5693_QOUT;
reg x_reg_L1_16__retimed_I5691_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5691_QOUT <= N9232;
	end
assign N10205 = x_reg_L1_16__retimed_I5691_QOUT;
reg x_reg_L1_15__retimed_I5689_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5689_QOUT <= N9227;
	end
assign N10200 = x_reg_L1_15__retimed_I5689_QOUT;
reg x_reg_L1_14__retimed_I5687_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5687_QOUT <= N9222;
	end
assign N10195 = x_reg_L1_14__retimed_I5687_QOUT;
reg x_reg_L1_13__retimed_I5685_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5685_QOUT <= N9217;
	end
assign N10190 = x_reg_L1_13__retimed_I5685_QOUT;
reg x_reg_L1_12__retimed_I5683_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5683_QOUT <= N9212;
	end
assign N10185 = x_reg_L1_12__retimed_I5683_QOUT;
reg x_reg_L1_11__retimed_I5681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5681_QOUT <= N9207;
	end
assign N10180 = x_reg_L1_11__retimed_I5681_QOUT;
reg x_reg_L1_10__retimed_I5679_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5679_QOUT <= N9202;
	end
assign N10175 = x_reg_L1_10__retimed_I5679_QOUT;
reg x_reg_L1_9__retimed_I5677_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5677_QOUT <= N9197;
	end
assign N10170 = x_reg_L1_9__retimed_I5677_QOUT;
reg x_reg_L1_8__retimed_I5675_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5675_QOUT <= N9192;
	end
assign N10165 = x_reg_L1_8__retimed_I5675_QOUT;
reg x_reg_L1_7__retimed_I5673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5673_QOUT <= N9187;
	end
assign N10160 = x_reg_L1_7__retimed_I5673_QOUT;
reg x_reg_L1_6__retimed_I5671_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5671_QOUT <= N9182;
	end
assign N10155 = x_reg_L1_6__retimed_I5671_QOUT;
reg x_reg_L1_5__retimed_I5669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5669_QOUT <= N9177;
	end
assign N10150 = x_reg_L1_5__retimed_I5669_QOUT;
reg x_reg_L1_4__retimed_I5667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5667_QOUT <= N9172;
	end
assign N10145 = x_reg_L1_4__retimed_I5667_QOUT;
reg x_reg_L1_3__retimed_I5665_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5665_QOUT <= N9167;
	end
assign N10140 = x_reg_L1_3__retimed_I5665_QOUT;
reg x_reg_L1_2__retimed_I5663_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5663_QOUT <= N9162;
	end
assign N10135 = x_reg_L1_2__retimed_I5663_QOUT;
reg x_reg_L1_1__retimed_I5661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5661_QOUT <= N9157;
	end
assign N10130 = x_reg_L1_1__retimed_I5661_QOUT;
reg x_reg_L1_0__retimed_I5659_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5659_QOUT <= N9152;
	end
assign N10125 = x_reg_L1_0__retimed_I5659_QOUT;
reg x_reg_L1_21__retimed_I5654_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5654_QOUT <= N9141;
	end
assign N10114 = x_reg_L1_21__retimed_I5654_QOUT;
reg x_reg_L1_20__retimed_I5650_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5650_QOUT <= N9132;
	end
assign N10105 = x_reg_L1_20__retimed_I5650_QOUT;
reg x_reg_L1_19__retimed_I5646_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5646_QOUT <= N9123;
	end
assign N10096 = x_reg_L1_19__retimed_I5646_QOUT;
reg x_reg_L1_18__retimed_I5642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5642_QOUT <= N9114;
	end
assign N10087 = x_reg_L1_18__retimed_I5642_QOUT;
reg x_reg_L1_17__retimed_I5638_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5638_QOUT <= N9105;
	end
assign N10078 = x_reg_L1_17__retimed_I5638_QOUT;
reg x_reg_L1_16__retimed_I5634_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5634_QOUT <= N9096;
	end
assign N10069 = x_reg_L1_16__retimed_I5634_QOUT;
reg x_reg_L1_15__retimed_I5630_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5630_QOUT <= N9087;
	end
assign N10060 = x_reg_L1_15__retimed_I5630_QOUT;
reg x_reg_L1_14__retimed_I5626_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5626_QOUT <= N9078;
	end
assign N10051 = x_reg_L1_14__retimed_I5626_QOUT;
reg x_reg_L1_13__retimed_I5622_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5622_QOUT <= N9069;
	end
assign N10042 = x_reg_L1_13__retimed_I5622_QOUT;
reg x_reg_L1_12__retimed_I5618_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5618_QOUT <= N9060;
	end
assign N10033 = x_reg_L1_12__retimed_I5618_QOUT;
reg x_reg_L1_11__retimed_I5614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5614_QOUT <= N9051;
	end
assign N10024 = x_reg_L1_11__retimed_I5614_QOUT;
reg x_reg_L1_10__retimed_I5610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5610_QOUT <= N9042;
	end
assign N10015 = x_reg_L1_10__retimed_I5610_QOUT;
reg x_reg_L1_9__retimed_I5606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5606_QOUT <= N9033;
	end
assign N10006 = x_reg_L1_9__retimed_I5606_QOUT;
reg x_reg_L1_8__retimed_I5602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5602_QOUT <= N9024;
	end
assign N9997 = x_reg_L1_8__retimed_I5602_QOUT;
reg x_reg_L1_7__retimed_I5598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5598_QOUT <= N9015;
	end
assign N9988 = x_reg_L1_7__retimed_I5598_QOUT;
reg x_reg_L1_6__retimed_I5594_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5594_QOUT <= N9006;
	end
assign N9979 = x_reg_L1_6__retimed_I5594_QOUT;
reg x_reg_L1_5__retimed_I5590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5590_QOUT <= N8997;
	end
assign N9970 = x_reg_L1_5__retimed_I5590_QOUT;
reg x_reg_L1_4__retimed_I5586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5586_QOUT <= N8988;
	end
assign N9961 = x_reg_L1_4__retimed_I5586_QOUT;
reg x_reg_L1_3__retimed_I5582_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5582_QOUT <= N8979;
	end
assign N9952 = x_reg_L1_3__retimed_I5582_QOUT;
reg x_reg_L1_2__retimed_I5578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5578_QOUT <= N8970;
	end
assign N9943 = x_reg_L1_2__retimed_I5578_QOUT;
reg x_reg_L1_1__retimed_I5574_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5574_QOUT <= N8961;
	end
assign N9934 = x_reg_L1_1__retimed_I5574_QOUT;
reg x_reg_L1_0__retimed_I5573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5573_QOUT <= N8958;
	end
assign N9931 = x_reg_L1_0__retimed_I5573_QOUT;
assign N13249 = !N9931;
assign N13250 = !N13249;
reg x_reg_L1_0__retimed_I5570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5570_QOUT <= N8952;
	end
assign N9925 = x_reg_L1_0__retimed_I5570_QOUT;
reg x_reg_L0_21__retimed_I5520_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5520_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26;
	end
assign N9758 = x_reg_L0_21__retimed_I5520_QOUT;
reg x_reg_L0_21__retimed_I5518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5518_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144;
	end
assign N9732 = x_reg_L0_21__retimed_I5518_QOUT;
reg x_reg_L0_21__retimed_I5516_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5516_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225;
	end
assign N9706 = x_reg_L0_21__retimed_I5516_QOUT;
reg x_reg_L1_22__retimed_I5514_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I5514_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053;
	end
assign N9680 = x_reg_L1_22__retimed_I5514_QOUT;
reg x_reg_L1_22__retimed_I5513_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I5513_QOUT <= N8945;
	end
assign N9678 = x_reg_L1_22__retimed_I5513_QOUT;
reg x_reg_L1_23__retimed_I5511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I5511_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004;
	end
assign N9673 = x_reg_L1_23__retimed_I5511_QOUT;
reg x_reg_L1_23__retimed_I5510_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I5510_QOUT <= N8938;
	end
assign N9671 = x_reg_L1_23__retimed_I5510_QOUT;
reg x_reg_L1_24__retimed_I5508_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I5508_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1];
	end
assign N9666 = x_reg_L1_24__retimed_I5508_QOUT;
reg x_reg_L1_25__retimed_I5505_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I5505_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2];
	end
assign N9659 = x_reg_L1_25__retimed_I5505_QOUT;
reg x_reg_L1_26__retimed_I5502_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I5502_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3];
	end
assign N9652 = x_reg_L1_26__retimed_I5502_QOUT;
reg x_reg_L1_27__retimed_I5499_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I5499_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4];
	end
assign N9645 = x_reg_L1_27__retimed_I5499_QOUT;
reg x_reg_L1_28__retimed_I5496_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I5496_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5];
	end
assign N9638 = x_reg_L1_28__retimed_I5496_QOUT;
reg x_reg_L1_29__retimed_I5494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I5494_QOUT <= N8900;
	end
assign N9633 = x_reg_L1_29__retimed_I5494_QOUT;
reg x_reg_L1_29__retimed_I5493_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I5493_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6];
	end
assign N9631 = x_reg_L1_29__retimed_I5493_QOUT;
reg x_reg_L1_30__retimed_I5490_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I5490_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7];
	end
assign N9624 = x_reg_L1_30__retimed_I5490_QOUT;
reg x_reg_L0_21__retimed_I5330_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5330_QOUT <= a_man[21];
	end
assign N9257 = x_reg_L0_21__retimed_I5330_QOUT;
reg x_reg_L0_20__retimed_I5328_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I5328_QOUT <= a_man[20];
	end
assign N9252 = x_reg_L0_20__retimed_I5328_QOUT;
reg x_reg_L0_19__retimed_I5326_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I5326_QOUT <= a_man[19];
	end
assign N9247 = x_reg_L0_19__retimed_I5326_QOUT;
reg x_reg_L0_18__retimed_I5324_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I5324_QOUT <= a_man[18];
	end
assign N9242 = x_reg_L0_18__retimed_I5324_QOUT;
reg x_reg_L0_17__retimed_I5322_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I5322_QOUT <= a_man[17];
	end
assign N9237 = x_reg_L0_17__retimed_I5322_QOUT;
reg x_reg_L0_16__retimed_I5320_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I5320_QOUT <= a_man[16];
	end
assign N9232 = x_reg_L0_16__retimed_I5320_QOUT;
reg x_reg_L0_15__retimed_I5318_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5318_QOUT <= a_man[15];
	end
assign N9227 = x_reg_L0_15__retimed_I5318_QOUT;
reg x_reg_L0_14__retimed_I5316_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I5316_QOUT <= a_man[14];
	end
assign N9222 = x_reg_L0_14__retimed_I5316_QOUT;
reg x_reg_L0_13__retimed_I5314_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I5314_QOUT <= a_man[13];
	end
assign N9217 = x_reg_L0_13__retimed_I5314_QOUT;
reg x_reg_L0_12__retimed_I5312_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I5312_QOUT <= a_man[12];
	end
assign N9212 = x_reg_L0_12__retimed_I5312_QOUT;
reg x_reg_L0_11__retimed_I5310_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I5310_QOUT <= a_man[11];
	end
assign N9207 = x_reg_L0_11__retimed_I5310_QOUT;
reg x_reg_L0_10__retimed_I5308_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I5308_QOUT <= a_man[10];
	end
assign N9202 = x_reg_L0_10__retimed_I5308_QOUT;
reg x_reg_L0_9__retimed_I5306_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I5306_QOUT <= a_man[9];
	end
assign N9197 = x_reg_L0_9__retimed_I5306_QOUT;
reg x_reg_L0_8__retimed_I5304_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I5304_QOUT <= a_man[8];
	end
assign N9192 = x_reg_L0_8__retimed_I5304_QOUT;
reg x_reg_L0_7__retimed_I5302_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I5302_QOUT <= a_man[7];
	end
assign N9187 = x_reg_L0_7__retimed_I5302_QOUT;
reg x_reg_L0_6__retimed_I5300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I5300_QOUT <= a_man[6];
	end
assign N9182 = x_reg_L0_6__retimed_I5300_QOUT;
reg x_reg_L0_5__retimed_I5298_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I5298_QOUT <= a_man[5];
	end
assign N9177 = x_reg_L0_5__retimed_I5298_QOUT;
reg x_reg_L0_4__retimed_I5296_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I5296_QOUT <= a_man[4];
	end
assign N9172 = x_reg_L0_4__retimed_I5296_QOUT;
reg x_reg_L0_3__retimed_I5294_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I5294_QOUT <= a_man[3];
	end
assign N9167 = x_reg_L0_3__retimed_I5294_QOUT;
reg x_reg_L0_2__retimed_I5292_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I5292_QOUT <= a_man[2];
	end
assign N9162 = x_reg_L0_2__retimed_I5292_QOUT;
reg x_reg_L0_1__retimed_I5290_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I5290_QOUT <= a_man[1];
	end
assign N9157 = x_reg_L0_1__retimed_I5290_QOUT;
reg x_reg_L0_0__retimed_I5288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5288_QOUT <= a_man[0];
	end
assign N9152 = x_reg_L0_0__retimed_I5288_QOUT;
reg x_reg_L0_21__retimed_I5283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5283_QOUT <= b_man[21];
	end
assign N9141 = x_reg_L0_21__retimed_I5283_QOUT;
reg x_reg_L0_20__retimed_I5279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I5279_QOUT <= b_man[20];
	end
assign N9132 = x_reg_L0_20__retimed_I5279_QOUT;
reg x_reg_L0_19__retimed_I5275_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I5275_QOUT <= b_man[19];
	end
assign N9123 = x_reg_L0_19__retimed_I5275_QOUT;
reg x_reg_L0_18__retimed_I5271_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I5271_QOUT <= b_man[18];
	end
assign N9114 = x_reg_L0_18__retimed_I5271_QOUT;
reg x_reg_L0_17__retimed_I5267_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I5267_QOUT <= b_man[17];
	end
assign N9105 = x_reg_L0_17__retimed_I5267_QOUT;
reg x_reg_L0_16__retimed_I5263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I5263_QOUT <= b_man[16];
	end
assign N9096 = x_reg_L0_16__retimed_I5263_QOUT;
reg x_reg_L0_15__retimed_I5259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5259_QOUT <= b_man[15];
	end
assign N9087 = x_reg_L0_15__retimed_I5259_QOUT;
reg x_reg_L0_14__retimed_I5255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I5255_QOUT <= b_man[14];
	end
assign N9078 = x_reg_L0_14__retimed_I5255_QOUT;
reg x_reg_L0_13__retimed_I5251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I5251_QOUT <= b_man[13];
	end
assign N9069 = x_reg_L0_13__retimed_I5251_QOUT;
reg x_reg_L0_12__retimed_I5247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I5247_QOUT <= b_man[12];
	end
assign N9060 = x_reg_L0_12__retimed_I5247_QOUT;
reg x_reg_L0_11__retimed_I5243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I5243_QOUT <= b_man[11];
	end
assign N9051 = x_reg_L0_11__retimed_I5243_QOUT;
reg x_reg_L0_10__retimed_I5239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I5239_QOUT <= b_man[10];
	end
assign N9042 = x_reg_L0_10__retimed_I5239_QOUT;
reg x_reg_L0_9__retimed_I5235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I5235_QOUT <= b_man[9];
	end
assign N9033 = x_reg_L0_9__retimed_I5235_QOUT;
reg x_reg_L0_8__retimed_I5231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I5231_QOUT <= b_man[8];
	end
assign N9024 = x_reg_L0_8__retimed_I5231_QOUT;
reg x_reg_L0_7__retimed_I5227_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I5227_QOUT <= b_man[7];
	end
assign N9015 = x_reg_L0_7__retimed_I5227_QOUT;
reg x_reg_L0_6__retimed_I5223_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I5223_QOUT <= b_man[6];
	end
assign N9006 = x_reg_L0_6__retimed_I5223_QOUT;
reg x_reg_L0_5__retimed_I5219_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I5219_QOUT <= b_man[5];
	end
assign N8997 = x_reg_L0_5__retimed_I5219_QOUT;
reg x_reg_L0_4__retimed_I5215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I5215_QOUT <= b_man[4];
	end
assign N8988 = x_reg_L0_4__retimed_I5215_QOUT;
reg x_reg_L0_3__retimed_I5211_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I5211_QOUT <= b_man[3];
	end
assign N8979 = x_reg_L0_3__retimed_I5211_QOUT;
reg x_reg_L0_2__retimed_I5207_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I5207_QOUT <= b_man[2];
	end
assign N8970 = x_reg_L0_2__retimed_I5207_QOUT;
reg x_reg_L0_1__retimed_I5203_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I5203_QOUT <= b_man[1];
	end
assign N8961 = x_reg_L0_1__retimed_I5203_QOUT;
reg x_reg_L0_0__retimed_I5202_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5202_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47;
	end
assign N8958 = x_reg_L0_0__retimed_I5202_QOUT;
reg x_reg_L0_0__retimed_I5199_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5199_QOUT <= b_man[0];
	end
assign N8952 = x_reg_L0_0__retimed_I5199_QOUT;
reg x_reg_L0_22__retimed_I5196_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5196_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055;
	end
assign N8945 = x_reg_L0_22__retimed_I5196_QOUT;
reg x_reg_L0_23__retimed_I5193_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I5193_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025;
	end
assign N8938 = x_reg_L0_23__retimed_I5193_QOUT;
reg x_reg_L0_29__retimed_I5177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_29__retimed_I5177_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008;
	end
assign N8900 = x_reg_L0_29__retimed_I5177_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007 = !(a_exp[0] & a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434 = !((a_exp[7] & a_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047 = !(((a_man[0] | a_man[1]) | a_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896 = !(b_exp[0] & b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426 = !((b_exp[7] & b_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936 = !(((b_man[0] | b_man[1]) | b_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919 = !(b_man[10] | b_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938 = !(b_man[6] | b_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927 = !(b_man[8] | b_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947 = !(b_man[4] | b_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092 = !(b_exp[0] | b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099 = !(b_exp[5] | b_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096 = !(b_exp[7] | b_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087 = !(b_exp[3] | b_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0] = (!b_exp[0]) ^ a_exp[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318 = (!b_man[22]) ^ b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217 = !a_man[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504 = !a_man[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862 = !a_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011 = b_man[22] | b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392 = (!b_man[20]) ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007 = b_man[21] ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552 = !b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415 = !a_man[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152 = !a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716 = !a_man[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076 = !a_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169 = b_man[19] ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463 = (!b_man[18]) ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407 = !b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529 = (!b_man[16]) ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973 = b_man[17] ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268 = !b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616 = !a_man[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352 = !a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924 = !a_man[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276 = !a_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212 = !a_man[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566 = !a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124 = !b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598 = (!b_man[14]) ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751 = b_man[15] ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664 = (!b_man[12]) ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942 = b_man[13] ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981 = !b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720 = b_man[11] ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737 = (!b_man[10]) ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827 = !b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131 = !a_man[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473 = !a_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417 = !a_man[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779 = !a_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805 = (!b_man[8]) ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911 = b_man[9] ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678 = !b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334 = !a_man[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675 = !a_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871 = (!b_man[6]) ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691 = b_man[7] ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531 = !b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881 = b_man[5] ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941 = (!b_man[4]) ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377 = !b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624 = !a_man[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988 = !a_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014 = (!b_man[2]) ^ b_man[1];
assign N13251 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014;
assign N13252 = !N13251;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662 = b_man[3] ^ b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237 = !b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357 & N13252) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268 = !a_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640 & N13252) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357 = !b_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721 = !(b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361 = !b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529 = !a_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831 = !(b_man[21] & b_man[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543 = !(b_man[19] & b_man[20]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901 = b_man[21] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610 = !(b_man[17] & b_man[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971 = b_man[19] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676 = !(b_man[15] & b_man[16]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043 = b_man[17] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749 = !(b_man[13] & b_man[14]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105 = b_man[15] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817 = !(b_man[11] & b_man[12]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172 = b_man[13] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883 = !(b_man[9] & b_man[10]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236 = b_man[11] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952 = !(b_man[7] & b_man[8]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301 = b_man[9] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028 = !(b_man[5] & b_man[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369 = b_man[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090 = !(b_man[3] & b_man[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430 = b_man[5] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154 = !(b_man[1] & b_man[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495 = b_man[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588) & (!N13252)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364) & (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678 = !(b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513) | (!(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739)));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107);
assign N13270 = !N11981;
assign N13273 = !(N11983 & N11829);
assign N13271 = !(N13270 & N13273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557 = !N13271;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557) & (!N11973)) | (!N11971);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440 = !(((N11962 & N11812) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441) | N11960);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707 = !(((N11664 | N11951) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440) & N11949);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707 & N11319) | N11941);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838;
assign N13280 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542 ^ N11930;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47] = !N13280;
assign N13319 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 = !N13319;
assign N13253 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360;
assign N13262 = !N13253;
assign N13261 = !N13253;
assign N13260 = !N13253;
assign N13259 = !N13253;
assign N13258 = !N13253;
assign N13257 = !N13253;
assign N13256 = !N13253;
assign N13255 = !N13253;
assign N13254 = !N13253;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707) ^ N11319;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[47] = !(N13254 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383 & N11343) | N11552);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336 ^ N11307;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440) & (!N11664)) | (!N11662);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914) ^ N11325;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44] = (N13256 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44]) | ((!N13256) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383) ^ N11343;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43] = (N13254 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43]) | ((!N13254) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914 & N11325) | N11539);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746 ^ N11301;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46] = (N13255 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46]) | ((!N13255) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45] = (N13255 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45]) | ((!N13255) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306 & N11684) | N11717);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176 ^ N11536;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163) & (!N11712)) | (!N11710);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325) ^ N11549;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36] = (N13257 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36]) | ((!N13257) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306) ^ N11684;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35] = (N13257 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35]) | ((!N13257) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325 & N11549) | N11573);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972 ^ N11337;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441 & N11812) | N11810);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643) ^ N11355;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38] = (N13256 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38]) | ((!N13256) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157 = !N12649;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497 = !N12652;
assign N13287 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235 = !N13287;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235 & N11906) | N11904);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522) & (!N11793)) | (!N11791);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376) ^ N11658;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34] = (N13258 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34]) | ((!N13258) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522 ^ N11672;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33] = (N13257 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33]) | ((!N13257) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958) & (!N11804)) | (!N11802);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879) ^ N11678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32] = (N13258 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32]) | ((!N13258) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958 ^ N11702;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31] = (N13257 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31]) | ((!N13257) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37] = (N13254 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37]) | ((!N13254) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595 & N11727) | N11742);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584 ^ N11583;
assign N13294 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557) & (!N11758)) | (!N11756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044 = !N13294;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044) ^ N11589;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28] = (N13257 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28]) | ((!N13257) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595) ^ N11727;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27] = (N13256 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27]) | ((!N13256) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044 & N11589) | N11592);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367 ^ N11361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30] = (N13256 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30]) | ((!N13256) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530 = !N12655;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886 = !N12658;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242 = !((N11829 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242) & (!N11823)) | (!N11821);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798) ^ N11733;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242 ^ N11739;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285 = !((N11829 & N11831) | N11840);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285 ^ N11752;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24] = (N13258 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24]) | ((!N13258) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29] = (N13255 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29]) | ((!N13255) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637) & (!N11694)) | (!N11692);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121 & N11349) | N11559);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550 ^ N11313;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42] = (N13255 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42]) | ((!N13255) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121) ^ N11349;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41] = (N13255 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41]) | ((!N13255) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643 & N11355) | N11566);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761 ^ N11331;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40] = (N13256 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40]) | ((!N13256) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39] = (N13254 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39]) | ((!N13254) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[24] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[47] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22] = (!N11829) ^ N11831;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[23] = (N13254 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23]) | ((!N13254) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23 = a_sign ^ b_sign;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[1] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[2] = (N13259 & N11467) | ((!N13259) & N11465);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[5] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[6] = (N13259 & N11488) | ((!N13259) & N11453);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[4] = (N13260 & N11451) | ((!N13260) & N11507);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[7] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[8] = (N13260 & N11472) | ((!N13260) & N11495);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[6]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[4]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[9] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[10] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[10] = (N13258 & N11460) | ((!N13258) & N11458);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[13] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[14] = (N13259 & N11481) | ((!N13259) & N11479);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[12] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[12] = (N13260 & N11502) | ((!N13260) & N11500);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[15] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[16] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[16] = (N13260 & N11523) | ((!N13260) & N11521);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[10] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[14]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[12]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[5] = (N13258 & N11453) | ((!N13258) & N11451);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[9] = (N13259 & N11458) | ((!N13259) & N11472);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[7] = (N13259 & N11495) | ((!N13259) & N11488);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[11] = (N13260 & N11500) | ((!N13260) & N11460);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[5] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[9]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[7]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[3] = (N13261 & N11507) | ((!N13261) & N11467);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21] = (!N11835) ^ N11837;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[22] = (N13262 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22]) | ((!N13262) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[3] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[20] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[20] = (N13261 & N12644) | ((!N13261) & N11624);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[17] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[18] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[18] = (N13262 & N11645) | ((!N13262) & N11643);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[20] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[0] = b_man[1] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[0] = N13261 & N11610;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[1] = (N13261 & N11465) | ((!N13261) & N11610);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[21] = (N13261 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21]) | ((!N13261) & N12644);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[13] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N11479) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N11502);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[17] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N11643) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N11523);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[15] = (N13262 & N11521) | ((!N13262) & N11481);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[19] = (N13262 & N11624) | ((!N13262) & N11645);
assign N13303 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[13] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[17]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[15]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[19]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679 = !N13303;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[1]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[21]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443) | N10969) | N10971) | N10973);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447 = ((N10921 | N10923) | N10925) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450 = ((!N10925) & (!N10923)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[23] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447);
assign N13309 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[24]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47]);
assign N13311 = !N13309;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 = !N13311;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10814) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10812);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765 = b_exp[0] | a_exp[0];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1]} = {1'B0, a_exp[1]} + {1'B0, b_exp[1]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0] | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1]));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2]} = {1'B0, a_exp[2]} + {1'B0, b_exp[2]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[2] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10860) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10858);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3]} = {1'B0, a_exp[3]} + {1'B0, b_exp[3]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4]} = {1'B0, a_exp[4]} + {1'B0, b_exp[4]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[4] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10869) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10867);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5]} = {1'B0, a_exp[5]} + {1'B0, b_exp[5]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10823) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10821);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6]} = {1'B0, a_exp[6]} + {1'B0, b_exp[6]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761 = !a_exp[7];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]} = {1'B0, b_exp[7]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10878) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10876);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10887) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10885);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8] = (!a_exp[7]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[8] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10800) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[6] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10832) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10830);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10841) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10839);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9] = !(a_exp[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N10792) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N10790);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964 = !(((N10751 | N10753) | N9758) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123 = !N12662;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 = !(N10567 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123);
assign N13263 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082;
assign N13264 = !N13263;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178 = !(N13264 & N10230);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[21] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 = N10645 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 = !(N10645 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10422) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10428));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 = !(N10593 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123);
assign N13265 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192;
assign N13266 = !N13265;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 = !(N10619 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123);
assign N13267 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106;
assign N13268 = !N13267;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986 = !(rm[0] & rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7 = !(rm[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173 = !((N13266 & N10114) | (N13268 & N13250));
assign x[21] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095 = !(N13264 & N10225);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[20] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10413) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10419));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199 = !((N13266 & N10105) | (N13268 & N13250));
assign x[20] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205 = !(N13264 & N10220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10404) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10410));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221 = !((N13266 & N10096) | (N13268 & N13250));
assign x[19] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120 = !(N13264 & N10215);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[18] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10395) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10401));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247 = !((N13266 & N10087) | (N13268 & N13250));
assign x[18] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228 = !(N13264 & N10210);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[17] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10386) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10392));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078 = !((N13266 & N10078) | (N13268 & N13250));
assign x[17] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146 = !(N13264 & N10205);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[16] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10377) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10383));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103 = !((N13266 & N10069) | (N13268 & N13250));
assign x[16] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061 = !(N13264 & N10200);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[15] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10368) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10374));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129 = !((N13266 & N10060) | (N13268 & N13250));
assign x[15] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168 = !(N13264 & N10195);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10359) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10365));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154 = !((N13266 & N10051) | (N13268 & N13250));
assign x[14] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085 = !(N13264 & N10190);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[13] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10350) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10356));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177 = !((N13266 & N10042) | (N13268 & N13250));
assign x[13] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193 = !(N13264 & N10185);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10341) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10347));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203 = !((N13266 & N10033) | (N13268 & N13250));
assign x[12] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110 = !(N13264 & N10180);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10332) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10338));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226 = !((N13266 & N10024) | (N13268 & N13250));
assign x[11] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216 = !(N13264 & N10175);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[10] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10323) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10329));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060 = !((N13266 & N10015) | (N13268 & N13250));
assign x[10] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135 = !(N13264 & N10170);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10314) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10320));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083 = !((N13266 & N10006) | (N13268 & N13250));
assign x[9] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242 = !(N13264 & N10165);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10305) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10311));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108 = !((N13266 & N9997) | (N13268 & N13250));
assign x[8] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162 = !(N13264 & N10160);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10296) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134 = !((N13266 & N9988) | (N13268 & N13250));
assign x[7] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073 = !(N13264 & N10155);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10287) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10293));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160 = !((N13266 & N9979) | (N13268 & N13250));
assign x[6] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185 = !(N13264 & N10150);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10278) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10284));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183 = !((N13266 & N9970) | (N13268 & N13250));
assign x[5] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100 = !(N13264 & N10145);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10269) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10275));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209 = !((N13266 & N9961) | (N13268 & N13250));
assign x[4] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210 = !(N13264 & N10140);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10260) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10266));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232 = !((N13266 & N9952) | (N13268 & N13250));
assign x[3] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126 = !(N13264 & N10135);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10251) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10257));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064 = !((N13266 & N9943) | (N13268 & N13250));
assign x[2] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234 = !(N13264 & N10130);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10242) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10248));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089 = !((N13266 & N9934) | (N13268 & N13250));
assign x[1] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150 = !(N13264 & N10125);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & N10233) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & N10239));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114 = !((N13266 & N9925) | (N13268 & N13250));
assign x[0] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[22]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47);
assign x[22] = !((N13248 & N9678) | ((!N13248) & N9680));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470;
assign x[30] = (N13248 & N9633) | ((!N13248) & N9624);
assign x[29] = (N13248 & N9633) | ((!N13248) & N9631);
assign x[28] = (N13248 & N9633) | ((!N13248) & N9638);
assign x[27] = (N13248 & N9633) | ((!N13248) & N9645);
assign x[26] = (N13248 & N9633) | ((!N13248) & N9652);
assign x[25] = (N13248 & N9633) | ((!N13248) & N9659);
assign x[24] = (N13248 & N9633) | ((!N13248) & N9666);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470);
assign x[23] = !((N13248 & N9671) | ((!N13248) & N9673));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22 & (!b_sign));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15 & a_sign) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23);
reg x_reg_L0_31__I1669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__I1669_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[31];
	end
assign N4120 = x_reg_L0_31__I1669_QOUT;
reg x_reg_L1_31__I1701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I1701_QOUT <= N4120;
	end
assign x[31] = x_reg_L1_31__I1701_QOUT;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  vbLxSAzaqhE= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



