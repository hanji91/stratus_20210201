/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:06:53 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_3 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__9,
	inst_cellmath__17;
wire [8:0] inst_cellmath__19;
wire [7:0] inst_cellmath__20;
wire [8:0] inst_cellmath__22;
wire  inst_cellmath__29,
	inst_cellmath__33,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42;
wire [18:0] inst_cellmath__51;
wire [24:0] inst_cellmath__60;
wire [39:0] inst_cellmath__62__W0, inst_cellmath__62__W1,
	inst_cellmath__63__W0, inst_cellmath__63__W1;
wire [39:0] inst_cellmath__64;
wire  inst_cellmath__67;
wire N447,N448,N449,N450,N451,N452,N453 
	,N454,N455,N456,N457,N477,N478,N479,N480 
	,N481,N482,N483,N484,N485,N486,N487,N488 
	,N489,N490,N491,N492,N493,N494,N495,N496 
	,N497,N498,N499,N500,N2353,N2355,N2376,N2378 
	,N2381,N2384,N2387,N2389,N2393,N2395,N2402,N2404 
	,N2408,N2444,N2449,N2451,N2454,N2457,N2459,N2464 
	,N2483,N2486,N2489,N2514,N2516,N2518,N2523,N2526 
	,N2576,N2577,N2578,N2579,N2580,N2581,N2583,N2584 
	,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592 
	,N2593,N2595,N2596,N2597,N2599,N2600,N2601,N2602 
	,N2603,N2604,N2605,N2606,N2608,N2609,N2610,N2611 
	,N2614,N2615,N2616,N2617,N2619,N2621,N2623,N2624 
	,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632 
	,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2641 
	,N2642,N2643,N2644,N2645,N2647,N2648,N2649,N2650 
	,N2652,N2655,N2656,N2658,N2659,N2660,N2661,N2663 
	,N2665,N2666,N2667,N2668,N2670,N2671,N2672,N2673 
	,N2674,N2675,N2677,N2678,N2679,N2680,N2681,N2682 
	,N2683,N2684,N2685,N2686,N2688,N2689,N2690,N2691 
	,N2694,N2695,N2696,N2697,N2698,N2699,N2701,N2702 
	,N2703,N2704,N2705,N2706,N2708,N2709,N2710,N2711 
	,N2712,N2713,N2714,N2715,N2717,N2719,N2720,N2721 
	,N2722,N2723,N2724,N2726,N2727,N2729,N2730,N2731 
	,N2732,N2734,N2735,N2736,N2738,N2739,N2741,N2742 
	,N2743,N2745,N2746,N2747,N2748,N2749,N2750,N2752 
	,N2753,N2754,N2755,N2758,N2760,N2762,N2763,N2764 
	,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773 
	,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2782 
	,N2783,N2784,N2785,N2787,N2788,N2789,N2790,N2791 
	,N2792,N2794,N2795,N2797,N2798,N2799,N2800,N2801 
	,N2802,N2803,N2804,N2806,N2809,N2810,N2811,N2812 
	,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820 
	,N2821,N2822,N2824,N2825,N2827,N2828,N2829,N2830 
	,N2831,N2832,N2833,N2834,N2835,N2837,N2838,N2839 
	,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848 
	,N2849,N2851,N2852,N2853,N2854,N2855,N2856,N2858 
	,N2859,N2861,N2862,N2863,N2865,N2866,N2868,N2869 
	,N2870,N2871,N2872,N2875,N2876,N2878,N2879,N2880 
	,N2881,N2882,N2884,N2885,N2886,N2887,N2888,N2889 
	,N2891,N2892,N2893,N2894,N2895,N2896,N3205,N3206 
	,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214 
	,N3215,N3216,N3218,N3219,N3220,N3221,N3222,N3223 
	,N3224,N3225,N3226,N3227,N3228,N3229,N3231,N3232 
	,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240 
	,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248 
	,N3249,N3250,N3252,N3253,N3254,N3255,N3256,N3257 
	,N3258,N3259,N3260,N3261,N3262,N3264,N3265,N3266 
	,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274 
	,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282 
	,N3283,N3284,N3285,N3287,N3288,N3289,N3290,N3291 
	,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299 
	,N3300,N3301,N3303,N3304,N3305,N3306,N3307,N3308 
	,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316 
	,N3317,N3318,N3319,N3320,N3322,N3323,N3324,N3325 
	,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333 
	,N3334,N3335,N3336,N3337,N3338,N3340,N3341,N3342 
	,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350 
	,N3351,N3352,N3354,N3355,N3356,N3357,N3358,N3359 
	,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367 
	,N3369,N3370,N3371,N3372,N3373,N3374,N3376,N3377 
	,N3378,N3379,N3380,N3381,N3382,N3383,N3384,N3385 
	,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394 
	,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402 
	,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410 
	,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418 
	,N3419,N3421,N3422,N3423,N3424,N3425,N3426,N3427 
	,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3436 
	,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444 
	,N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452 
	,N3453,N3454,N3455,N3457,N3458,N3459,N3460,N3461 
	,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469 
	,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478 
	,N3479,N3480,N3481,N3482,N3483,N3485,N3486,N3487 
	,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496 
	,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504 
	,N3505,N3506,N3507,N3508,N3510,N3511,N3512,N3513 
	,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521 
	,N3522,N3523,N3524,N3525,N3526,N3528,N3529,N3530 
	,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538 
	,N3539,N3540,N3541,N3542,N3543,N3545,N3546,N3547 
	,N3548,N3549,N3550,N3551,N3552,N3553,N3555,N3556 
	,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564 
	,N3565,N3566,N3567,N3568,N3569,N3570,N3571,N3572 
	,N3573,N3574,N3576,N3577,N3578,N3579,N3580,N3581 
	,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589 
	,N3590,N3592,N3593,N3594,N3595,N3596,N3597,N3598 
	,N3599,N3600,N3601,N3602,N3603,N3605,N3606,N3607 
	,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3616 
	,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624 
	,N3625,N3626,N3627,N3628,N3629,N3631,N3632,N3633 
	,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641 
	,N3642,N3643,N3645,N3646,N3647,N3648,N3649,N3650 
	,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658 
	,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3668 
	,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676 
	,N3677,N3679,N3680,N3681,N3682,N3683,N3684,N3685 
	,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693 
	,N3694,N3695,N3696,N3697,N3699,N3700,N3701,N3702 
	,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710 
	,N3711,N3713,N3714,N3715,N3716,N3717,N3718,N3719 
	,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727 
	,N3728,N3729,N3731,N3732,N3733,N3734,N3735,N3736 
	,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744 
	,N3745,N3746,N3748,N3749,N3750,N3751,N3752,N3753 
	,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761 
	,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770 
	,N3771,N3772,N3773,N3775,N3776,N3777,N3778,N3779 
	,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788 
	,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796 
	,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805 
	,N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813 
	,N3814,N3815,N3816,N3818,N3819,N3820,N3821,N3822 
	,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830 
	,N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839 
	,N3840,N3841,N3842,N3844,N3845,N3846,N3847,N3848 
	,N3849,N3850,N3852,N3853,N3854,N3855,N3856,N3857 
	,N3858,N3859,N3860,N3861,N3862,N3863,N3864,N3866 
	,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874 
	,N3875,N3876,N3878,N3879,N3880,N3881,N3882,N3883 
	,N3884,N3885,N3886,N3887,N3888,N3889,N3891,N3892 
	,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3901 
	,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909 
	,N3910,N3911,N3912,N3913,N3914,N3915,N3917,N3918 
	,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926 
	,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3935 
	,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943 
	,N3944,N3945,N3946,N3947,N3948,N3949,N3951,N3952 
	,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960 
	,N3961,N3964,N3965,N3966,N3967,N3968,N3969,N3970 
	,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978 
	,N3979,N3981,N3982,N3983,N3984,N3985,N3986,N3987 
	,N3988,N3989,N3990,N3991,N3992,N3994,N3995,N3996 
	,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004 
	,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013 
	,N4014,N4015,N4017,N4018,N4019,N4020,N4021,N4022 
	,N4023,N4024,N4025,N4026,N4027,N4029,N4030,N4031 
	,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039 
	,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4048 
	,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056 
	,N4057,N4058,N4059,N4061,N4062,N4063,N4064,N4065 
	,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074 
	,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082 
	,N4084,N4085,N4086,N4087,N4088,N4089,N4090,N4091 
	,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099 
	,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4108 
	,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116 
	,N4117,N4118,N4119,N4120,N4122,N4123,N4124,N4125 
	,N4126,N4127,N4128,N4129,N4130,N4132,N4133,N4134 
	,N4135,N4136,N4137,N5064,N5066,N5068,N5069,N5071 
	,N5072,N5073,N5074,N5075,N5077,N5078,N5079,N5080 
	,N5081,N5082,N5083,N5085,N5086,N5087,N5088,N5089 
	,N5090,N5091,N5092,N5093,N5094,N5096,N5097,N5099 
	,N5100,N5101,N5104,N5106,N5107,N5108,N5110,N5112 
	,N5113,N5114,N5115,N5116,N5117,N5118,N5120,N5121 
	,N5122,N5123,N5124,N5125,N5127,N5128,N5129,N5131 
	,N5132,N5133,N5134,N5135,N5136,N5137,N5139,N5140 
	,N5141,N5143,N5145,N5146,N5147,N5148,N5149,N5150 
	,N5152,N5153,N5154,N5155,N5156,N5157,N5158,N5159 
	,N5160,N5163,N5164,N5165,N5166,N5167,N5168,N5169 
	,N5171,N5173,N5174,N5175,N5176,N5177,N5178,N5179 
	,N5180,N5181,N5184,N5185,N5186,N5187,N5188,N5189 
	,N5191,N5192,N5194,N5195,N5196,N5197,N5198,N5199 
	,N5200,N5201,N5203,N5205,N5206,N5207,N5208,N5209 
	,N5210,N5211,N5213,N5214,N5216,N5217,N5218,N5219 
	,N5220,N5221,N5222,N5223,N5225,N5226,N5228,N5230 
	,N5231,N5233,N5234,N5235,N5236,N5237,N5238,N5239 
	,N5240,N5242,N5243,N5244,N5246,N5247,N5248,N5249 
	,N5250,N5251,N5252,N5254,N5256,N5257,N5258,N5259 
	,N5260,N5261,N5262,N5263,N5265,N5266,N5267,N5268 
	,N5269,N5270,N5271,N5272,N5274,N5275,N5276,N5278 
	,N5279,N5280,N5281,N5282,N5283,N5285,N5286,N5288 
	,N5289,N5291,N5292,N5293,N5294,N5295,N5297,N5298 
	,N5299,N5301,N5302,N5303,N5304,N5305,N5306,N5307 
	,N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5317 
	,N5318,N5320,N5321,N5322,N5323,N5324,N5325,N5326 
	,N5327,N5328,N5329,N5330,N5332,N5334,N5335,N5336 
	,N5337,N5339,N5340,N5341,N5342,N5343,N5344,N5345 
	,N5346,N5347,N5348,N5349,N5351,N5354,N5355,N5356 
	,N5357,N5358,N5359,N5360,N5363,N5364,N5365,N5366 
	,N5367,N5368,N5369,N5370,N5372,N5373,N5374,N5376 
	,N5378,N5379,N5380,N5381,N5382,N5383,N5384,N5386 
	,N5387,N5388,N5389,N5390,N5391,N5392,N5393,N5395 
	,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5723 
	,N5724,N5725,N5726,N5728,N5730,N5731,N5732,N5733 
	,N5734,N5735,N5736,N5737,N5738,N5739,N5740,N5741 
	,N5742,N5743,N5744,N5745,N5746,N5747,N5749,N5750 
	,N5751,N5753,N5754,N5755,N5756,N5758,N5759,N5760 
	,N5761,N5762,N5764,N5765,N5766,N5767,N5768,N5769 
	,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778 
	,N5779,N5780,N5781,N5782,N5784,N5785,N5786,N5787 
	,N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5797 
	,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5806 
	,N5807,N5808,N5809,N5810,N5811,N5812,N5813,N5814 
	,N5815,N5816,N5818,N5820,N5821,N5822,N5823,N5824 
	,N5825,N5826,N5827,N5829,N5830,N5831,N5833,N5834 
	,N5835,N5836,N5838,N5839,N5840,N5841,N5842,N5843 
	,N5844,N5846,N5847,N5848,N5849,N5850,N5851,N5852 
	,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860 
	,N5861,N5863,N5864,N5865,N5866,N5867,N5869,N5870 
	,N5872,N5873,N5874,N5875,N5876,N5877,N5879,N5880 
	,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888 
	,N5889,N5890,N5891,N5892,N5894,N5895,N5896,N5897 
	,N5898,N5899,N5900,N5901,N5903,N5904,N5905,N5906 
	,N5907,N5908,N5911,N5912,N5914,N5915,N5916,N5917 
	,N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5927 
	,N5928,N5929,N5930,N5931,N5932,N5933,N5934,N5935 
	,N5937,N5938,N5939,N5940,N5941,N5943,N5944,N5946 
	,N5947,N5948,N5949,N5950,N5951,N5952,N5954,N5955 
	,N5956,N5957,N5958,N5960,N5961,N5962,N5963,N5964 
	,N5965,N5966,N5967,N5968,N5969,N5970,N5971,N5972 
	,N5973,N5975,N5976,N5977,N5978,N5979,N5980,N5981 
	,N5982,N5983,N5984,N5985,N5986,N5987,N5988,N5989 
	,N5990,N5992,N5993,N5994,N5995,N5996,N5997,N5998 
	,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6007 
	,N6009,N6010,N6011,N6012,N6013,N6014,N6016,N6017 
	,N6018,N6019,N6021,N6022,N6023,N6024,N6026,N6027 
	,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035 
	,N6036,N6037,N6038,N6039,N6040,N6041,N6042,N6043 
	,N6046,N6047,N6048,N6049,N6051,N6052,N6053,N6055 
	,N6056,N6057,N6058,N6060,N6061,N6062,N6063,N6064 
	,N6065,N6066,N6067,N6069,N6070,N6071,N6072,N6073 
	,N6074,N6075,N6076,N6077,N6078,N6079,N6080,N6081 
	,N6082,N6084,N6085,N6086,N6087,N6088,N6089,N6091 
	,N6092,N6093,N6095,N6096,N6097,N6098,N6100,N6101 
	,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6109 
	,N6111,N6112,N6115,N6116,N6117,N6118,N6119,N6120 
	,N6121,N6122,N6123,N6124,N6126,N6127,N6128,N6130 
	,N6131,N6132,N6133,N6134,N6136,N6137,N6138,N6139 
	,N6140,N6141,N6142,N6143,N6145,N6146,N6147,N6148 
	,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156 
	,N6157,N6158,N6160,N6161,N6162,N6163,N6164,N6165 
	,N6167,N6168,N6169,N6170,N6171,N6172,N6173,N6174 
	,N6176,N6177,N6179,N6180,N6181,N6182,N6183,N6184 
	,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192 
	,N6194,N6195,N6196,N6197,N6198,N6199,N6200,N6201 
	,N6203,N6204,N6205,N6206,N6208,N6209,N6211,N6212 
	,N6213,N6214,N6215,N6216,N6217,N6218,N6219,N6220 
	,N6222,N6223,N6224,N6225,N6226,N6227,N6228,N6229 
	,N6230,N6232,N6233,N6234,N6235,N6236,N6239,N6240 
	,N6242,N6243,N6244,N6245,N6246,N6247,N6248,N6249 
	,N6250,N6251,N6252,N6253,N6255,N6256,N6257,N6258 
	,N6259,N6260,N6261,N6262,N6263,N6264,N6265,N6266 
	,N6267,N6268,N6269,N6270,N6272,N6273,N6275,N6276 
	,N6277,N6278,N6280,N6281,N6282,N6283,N6284,N6285 
	,N6286,N6287,N6289,N6290,N6291,N6292,N6293,N6294 
	,N6295,N6296,N6297,N6298,N6299,N6301,N6302,N6303 
	,N6304,N6305,N6306,N6307,N6308,N6309,N6310,N6311 
	,N6312,N6315,N6316,N6317,N6318,N6320,N6321,N6322 
	,N6324,N6325,N6326,N6327,N6328,N6329,N6331,N6332 
	,N6333,N6334,N6335,N6337,N6338,N6339,N6340,N6341 
	,N6342,N6343,N6344,N6345,N6346,N6347,N6348,N6349 
	,N6350,N6352,N6353,N6354,N6356,N6357,N6358,N6359 
	,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367 
	,N6369,N6370,N6371,N6372,N6373,N6374,N6375,N6376 
	,N6377,N6378,N6379,N6380,N6382,N6383,N6384,N6386 
	,N6387,N6388,N6389,N6390,N6391,N6392,N6393,N6394 
	,N6396,N6397,N6398,N6400,N6401,N6403,N6404,N6405 
	,N6406,N6407,N6408,N6409,N6410,N6412,N6413,N6414 
	,N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422 
	,N6424,N6425,N6427,N6428,N6429,N6430,N6432,N6433 
	,N6434,N6435,N6436,N6437,N6438,N6439,N6441,N6442 
	,N6444,N6445,N6446,N6447,N6448,N6449,N6450,N6451 
	,N6452,N6453,N6454,N6455,N6456,N6457,N6458,N6459 
	,N6461,N6462,N6463,N6464,N6465,N6467,N6468,N6469 
	,N6471,N6472,N6473,N6474,N6475,N6476,N6477,N6479 
	,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487 
	,N6488,N6489,N6490,N6492,N6493,N6494,N6495,N6496 
	,N6497,N6498,N6500,N6501,N6502,N6503,N6504,N6505 
	,N6508,N6509,N6511,N6512,N6513,N6514,N6515,N6516 
	,N6517,N6518,N6519,N6521,N6522,N6523,N6524,N6525 
	,N6526,N6527,N6528,N6529,N6530,N6531,N6532,N6533 
	,N6534,N6535,N6536,N6537,N6538,N6539,N6540,N6542 
	,N6543,N6545,N6546,N6547,N6548,N6549,N6550,N6551 
	,N6552,N6553,N6554,N6555,N6557,N6558,N6559,N6560 
	,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568 
	,N6570,N6571,N6572,N6574,N6575,N6576,N6577,N6578 
	,N6579,N6580,N6581,N7410,N7415,N7417,N7418,N7419 
	,N7420,N7425,N7427,N7429,N7430,N7434,N7437,N7439 
	,N7442,N7444,N7447,N7450,N7451,N7452,N7457,N7459 
	,N7460,N7462,N7464,N7465,N7468,N7471,N7474,N7476 
	,N7478,N7481,N7484,N7486,N7487,N7488,N7489,N7491 
	,N7492,N7497,N7499,N7500,N7501,N7503,N7508,N7511 
	,N7514,N7515,N7520,N7521,N7523,N7524,N7530,N7532 
	,N7533,N7535,N7540,N7542,N7543,N7545,N7546,N7550 
	,N7552,N7553,N7557,N7558,N7561,N7562,N7563,N7564 
	,N7565,N7567,N7568,N7570,N7571,N7572,N7575,N7578 
	,N7579,N7580,N7582,N7583,N7585,N7586,N7588,N7589 
	,N7590,N7592,N7593,N7597,N7599,N7601,N7605,N7606 
	,N7608,N7610,N7612,N7614,N7615,N7618,N7620,N7622 
	,N7623,N7627,N7629,N7631,N7634,N7635,N7638,N7640 
	,N7643,N7645,N7646,N7648,N7649,N7651,N7653,N7654 
	,N7655,N7659,N7663,N7664,N7667,N7668,N7670,N7674 
	,N7675,N7677,N7679,N7683,N7686,N7690,N7699,N7700 
	,N7702,N7703,N7704,N7706,N7709,N7712,N7716,N7719 
	,N7721,N7722,N7724,N7725,N7728,N7730,N7732,N7733 
	,N7735,N7736,N7741,N7744,N7745,N7747,N7748,N7749 
	,N7750,N7753,N7754,N7756,N7757,N7758,N7761,N7763 
	,N7767,N7769,N7770,N7771,N7772,N7776,N7777,N7778 
	,N7780,N7781,N7782,N7783,N7784,N7787,N7789,N7791 
	,N7794,N7795,N7797,N7798,N7799,N7800,N7802,N7803 
	,N7806,N7807,N7809,N7811,N7813,N7817,N7820,N7821 
	,N7823,N7824,N7826,N7829,N7831,N7832,N7834,N7837 
	,N7838,N7840,N7841,N7844,N7847,N7849,N7851,N7853 
	,N7856,N7857,N7858,N7861,N7862,N7864,N7866,N7868 
	,N7869,N7874,N7875,N7876,N7880,N7884,N7886,N7888 
	,N7890,N7892,N7894,N7895,N7896,N7899,N7902,N7904 
	,N7906,N7909,N7911,N7914,N7916,N7917,N7919,N7924 
	,N7926,N7927,N7929,N7936,N7937,N7939,N7940,N7941 
	,N7942,N7945,N7947,N7948,N7952,N7957,N7960,N7961 
	,N7963,N7964,N7965,N7968,N7969,N7971,N7972,N7973 
	,N7976,N7979,N7980,N7982,N7983,N7984,N7985,N7988 
	,N7989,N7991,N7992,N7995,N7996,N7998,N8001,N8003 
	,N8005,N8006,N8009,N8010,N8012,N8013,N8016,N8017 
	,N8018,N8022,N8024,N11653,N11660,N11661,N11662,N11669 
	,N11670,N11688,N11689,N11693,N11697,N11706,N11708,N11719 
	,N11728,N11739,N11743,N11749,N11756,N11758,N11788,N11795 
	;
NAND2XL inst_cellmath__9_0_I160 (.Y(N2353), .A(a_exp[7]), .B(a_exp[0]));
AND4XL inst_cellmath__9_0_I14164 (.Y(N2355), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL hyperpropagate_4_1_A_I5089 (.Y(N11743), .A(a_exp[6]), .B(a_exp[5]), .C(N2355));
NOR2XL hyperpropagate_4_1_A_I5090 (.Y(inst_cellmath__9), .A(N2353), .B(N11743));
NOR2XL inst_cellmath__15__5__I169 (.Y(N2381), .A(a_man[18]), .B(a_man[17]));
NOR2XL inst_cellmath__15__5__I173 (.Y(N2376), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__15__5__I174 (.Y(N2384), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__15__5__I175 (.Y(N2395), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__15__5__I176 (.Y(N2404), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__15__5__I14165 (.Y(N2389), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__15__5__I14166 (.Y(N2408), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 inst_cellmath__15__5__I14167 (.Y(N2402), .AN(N2381), .B(a_man[16]), .C(N2408), .D(a_man[15]));
NOR4X1 inst_cellmath__15__5__I180 (.Y(N2393), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N2389));
NAND4XL inst_cellmath__15__5__I182 (.Y(N2387), .A(N2376), .B(N2395), .C(N2384), .D(N2404));
NAND2XL inst_cellmath__15__5__I183 (.Y(N2378), .A(N2393), .B(N2402));
NOR2XL inst_cellmath__15__5__I184 (.Y(inst_cellmath__19[0]), .A(N2387), .B(N2378));
NOR2BX1 cynw_cm_float_rcp_I185 (.Y(inst_cellmath__29), .AN(inst_cellmath__9), .B(inst_cellmath__19[0]));
NOR2BX1 cynw_cm_float_rcp_I186 (.Y(x[31]), .AN(a_sign), .B(inst_cellmath__29));
INVXL cynw_cm_float_rcp_I5 (.Y(inst_cellmath__20[0]), .A(a_exp[0]));
INVXL cynw_cm_float_rcp_I6 (.Y(inst_cellmath__20[1]), .A(a_exp[1]));
INVXL cynw_cm_float_rcp_I8 (.Y(inst_cellmath__20[3]), .A(a_exp[3]));
INVXL cynw_cm_float_rcp_I10 (.Y(inst_cellmath__20[5]), .A(a_exp[5]));
INVXL cynw_cm_float_rcp_I12 (.Y(inst_cellmath__20[7]), .A(a_exp[7]));
ADDHX1 inst_cellmath__22_0_I188 (.CO(N2464), .S(inst_cellmath__22[0]), .A(inst_cellmath__20[0]), .B(inst_cellmath__19[0]));
XNOR2X1 inst_cellmath__22_0_I189 (.Y(inst_cellmath__22[1]), .A(inst_cellmath__20[1]), .B(N2464));
NOR2XL inst_cellmath__22_0_I190 (.Y(N2459), .A(inst_cellmath__20[1]), .B(N2464));
XNOR2X1 inst_cellmath__22_0_I191 (.Y(inst_cellmath__22[2]), .A(a_exp[2]), .B(N2459));
NAND2XL inst_cellmath__22_0_I192 (.Y(N2457), .A(a_exp[2]), .B(N2459));
XNOR2X1 inst_cellmath__22_0_I193 (.Y(inst_cellmath__22[3]), .A(inst_cellmath__20[3]), .B(N2457));
NOR2XL inst_cellmath__22_0_I194 (.Y(N2454), .A(inst_cellmath__20[3]), .B(N2457));
XNOR2X1 inst_cellmath__22_0_I195 (.Y(inst_cellmath__22[4]), .A(a_exp[4]), .B(N2454));
NAND2XL inst_cellmath__22_0_I196 (.Y(N2451), .A(a_exp[4]), .B(N2454));
XNOR2X1 inst_cellmath__22_0_I197 (.Y(inst_cellmath__22[5]), .A(inst_cellmath__20[5]), .B(N2451));
NOR2XL inst_cellmath__22_0_I198 (.Y(N2449), .A(inst_cellmath__20[5]), .B(N2451));
XNOR2X1 inst_cellmath__22_0_I199 (.Y(inst_cellmath__22[6]), .A(a_exp[6]), .B(N2449));
NAND2XL inst_cellmath__22_0_I200 (.Y(N2444), .A(a_exp[6]), .B(N2449));
XNOR2X1 inst_cellmath__22_0_I201 (.Y(inst_cellmath__22[7]), .A(inst_cellmath__20[7]), .B(N2444));
NOR2XL inst_cellmath__22_0_I202 (.Y(inst_cellmath__22[8]), .A(inst_cellmath__20[7]), .B(N2444));
NOR3XL inst_cellmath__17__6__I203 (.Y(N2486), .A(inst_cellmath__22[2]), .B(inst_cellmath__22[3]), .C(inst_cellmath__22[5]));
NOR2XL inst_cellmath__17__6__I204 (.Y(N2489), .A(inst_cellmath__22[6]), .B(inst_cellmath__22[7]));
NOR4BX1 inst_cellmath__17__6__I205 (.Y(N2483), .AN(N2489), .B(inst_cellmath__22[0]), .C(inst_cellmath__22[4]), .D(inst_cellmath__22[1]));
AO21XL cynw_cm_float_rcp_I5038 (.Y(inst_cellmath__17), .A0(N2486), .A1(N2483), .B0(inst_cellmath__22[8]));
MX2XL cynw_cm_float_rcp_I5073 (.Y(N447), .A(inst_cellmath__17), .B(inst_cellmath__19[0]), .S0(inst_cellmath__9));
NOR2BX1 cynw_cm_float_rcp_I210 (.Y(inst_cellmath__33), .AN(N447), .B(inst_cellmath__29));
NOR2XL inst_cellmath__34_0_I211 (.Y(N2523), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL inst_cellmath__34_0_I212 (.Y(N2526), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL inst_cellmath__34_0_I213 (.Y(N2514), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL inst_cellmath__34_0_I214 (.Y(N2518), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL inst_cellmath__34_0_I215 (.Y(N2516), .A(N2523), .B(N2514), .C(N2526), .D(N2518));
NOR2XL inst_cellmath__34_0_I216 (.Y(inst_cellmath__34), .A(N2516), .B(inst_cellmath__29));
NOR3XL cynw_cm_float_rcp_I217 (.Y(inst_cellmath__42), .A(inst_cellmath__29), .B(inst_cellmath__34), .C(inst_cellmath__33));
OR2XL cynw_cm_float_rcp_I218 (.Y(inst_cellmath__38), .A(inst_cellmath__29), .B(inst_cellmath__34));
MX2XL inst_cellmath__43_0_I219 (.Y(x[23]), .A(inst_cellmath__38), .B(inst_cellmath__22[0]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I220 (.Y(x[24]), .A(inst_cellmath__38), .B(inst_cellmath__22[1]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I221 (.Y(x[25]), .A(inst_cellmath__38), .B(inst_cellmath__22[2]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I222 (.Y(x[26]), .A(inst_cellmath__38), .B(inst_cellmath__22[3]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I223 (.Y(x[27]), .A(inst_cellmath__38), .B(inst_cellmath__22[4]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I224 (.Y(x[28]), .A(inst_cellmath__38), .B(inst_cellmath__22[5]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I225 (.Y(x[29]), .A(inst_cellmath__38), .B(inst_cellmath__22[6]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I226 (.Y(x[30]), .A(inst_cellmath__38), .B(inst_cellmath__22[7]), .S0(inst_cellmath__42));
OR4X1 cynw_cm_float_rcp_I227 (.Y(N448), .A(inst_cellmath__19[0]), .B(inst_cellmath__29), .C(inst_cellmath__34), .D(inst_cellmath__33));
INVXL cynw_cm_float_rcp_I24 (.Y(inst_cellmath__67), .A(N448));
INVXL cynw_cm_float_rcp_I25 (.Y(inst_cellmath__63__W0[33]), .A(a_man[15]));
INVX1 inst_cellmath__60_0_I228 (.Y(N2631), .A(a_man[4]));
INVXL inst_cellmath__60_0_I4950 (.Y(N11653), .A(N2631));
INVXL inst_cellmath__60_0_I4958 (.Y(N11661), .A(N11653));
INVX2 inst_cellmath__60_0_I4957 (.Y(N11660), .A(N11653));
INVXL inst_cellmath__60_0_I229 (.Y(N2698), .A(a_man[5]));
INVX1 inst_cellmath__60_0_I4959 (.Y(N11662), .A(N2698));
INVXL inst_cellmath__60_0_I4967 (.Y(N11670), .A(N11662));
INVX2 inst_cellmath__60_0_I4966 (.Y(N11669), .A(N11662));
INVX2 inst_cellmath__60_0_I230 (.Y(N2773), .A(a_man[6]));
INVXL inst_cellmath__60_0_I231 (.Y(N2579), .A(a_man[7]));
BUFX3 inst_cellmath__60_0_I5041 (.Y(N11688), .A(N2579));
INVXL inst_cellmath__60_0_I232 (.Y(N2648), .A(a_man[8]));
INVXL inst_cellmath__60_0_I4986 (.Y(N11689), .A(N2648));
INVX1 inst_cellmath__60_0_I4994 (.Y(N11697), .A(N11689));
INVXL inst_cellmath__60_0_I4990 (.Y(N11693), .A(N11689));
INVXL inst_cellmath__60_0_I233 (.Y(N2747), .A(a_man[9]));
BUFX2 inst_cellmath__60_0_I5042 (.Y(N11706), .A(N2747));
INVX2 inst_cellmath__60_0_I5005 (.Y(N11708), .A(a_man[10]));
INVXL inst_cellmath__60_0_I235 (.Y(N2888), .A(a_man[11]));
BUFX2 inst_cellmath__60_0_I5043 (.Y(N11719), .A(N2888));
INVXL inst_cellmath__60_0_I236 (.Y(N2637), .A(a_man[12]));
BUFX2 inst_cellmath__60_0_I5044 (.Y(N11728), .A(N2637));
INVX1 inst_cellmath__60_0_I237 (.Y(N2705), .A(a_man[13]));
INVXL inst_cellmath__60_0_I238 (.Y(N2777), .A(a_man[14]));
INVXL inst_cellmath__60_0_I239 (.Y(N2848), .A(inst_cellmath__63__W0[33]));
INVX2 inst_cellmath__60_0_I240 (.Y(N2876), .A(a_man[3]));
NOR2XL inst_cellmath__60_0_I244 (.Y(N2675), .A(N2876), .B(N2773));
NOR2XL inst_cellmath__60_0_I245 (.Y(N2822), .A(N2876), .B(N2579));
NOR2XL inst_cellmath__60_0_I246 (.Y(N2636), .A(N2876), .B(N11697));
NOR2XL inst_cellmath__60_0_I247 (.Y(N2779), .A(N2876), .B(N11706));
NOR2XL inst_cellmath__60_0_I248 (.Y(N2595), .A(N2876), .B(N11708));
NOR2XL inst_cellmath__60_0_I249 (.Y(N2732), .A(N2876), .B(N2888));
NOR2XL inst_cellmath__60_0_I250 (.Y(N2878), .A(N2876), .B(N2637));
NOR2XL inst_cellmath__60_0_I251 (.Y(N2691), .A(N2876), .B(N2705));
NOR2XL inst_cellmath__60_0_I252 (.Y(N2839), .A(N2876), .B(N2777));
OR2XL inst_cellmath__60_0_I253 (.Y(N2611), .A(N2876), .B(N2848));
NOR2XL inst_cellmath__60_0_I254 (.Y(N2815), .A(N11661), .B(N11670));
NOR2XL inst_cellmath__60_0_I255 (.Y(N2629), .A(N2631), .B(N2773));
NOR2XL inst_cellmath__60_0_I256 (.Y(N2771), .A(N11660), .B(N11688));
NOR2XL inst_cellmath__60_0_I257 (.Y(N2590), .A(N11660), .B(N11697));
NOR2XL inst_cellmath__60_0_I258 (.Y(N2727), .A(N2631), .B(N2747));
NOR2XL inst_cellmath__60_0_I259 (.Y(N2868), .A(N11660), .B(N11708));
NOR2XL inst_cellmath__60_0_I260 (.Y(N2685), .A(N11660), .B(N11719));
NOR2XL inst_cellmath__60_0_I261 (.Y(N2834), .A(N11661), .B(N11728));
NOR2XL inst_cellmath__60_0_I262 (.Y(N2647), .A(N11661), .B(N2705));
NOR2XL inst_cellmath__60_0_I263 (.Y(N2790), .A(N11661), .B(N2777));
OR2XL inst_cellmath__60_0_I264 (.Y(N2679), .A(N11661), .B(N2848));
NOR2XL inst_cellmath__60_0_I266 (.Y(N2763), .A(N11669), .B(N2773));
NOR2XL inst_cellmath__60_0_I267 (.Y(N2585), .A(N11669), .B(N11688));
NOR2XL inst_cellmath__60_0_I268 (.Y(N2721), .A(N2698), .B(N2648));
NOR2XL inst_cellmath__60_0_I269 (.Y(N2862), .A(N11669), .B(N11706));
NOR2XL inst_cellmath__60_0_I270 (.Y(N2680), .A(N11669), .B(N11708));
NOR2XL inst_cellmath__60_0_I271 (.Y(N2830), .A(N11670), .B(N11719));
NOR2XL inst_cellmath__60_0_I272 (.Y(N2643), .A(N11670), .B(N11728));
NOR2XL inst_cellmath__60_0_I273 (.Y(N2785), .A(N11670), .B(N2705));
NOR2XL inst_cellmath__60_0_I274 (.Y(N2602), .A(N11670), .B(N2777));
OR2XL inst_cellmath__60_0_I275 (.Y(N2753), .A(N11669), .B(N2848));
INVXL inst_cellmath__60_0_I276 (.Y(N2616), .A(N2773));
NOR2XL inst_cellmath__60_0_I277 (.Y(N2578), .A(N2773), .B(N11688));
NOR2XL inst_cellmath__60_0_I278 (.Y(N2715), .A(N2773), .B(N11697));
NOR2XL inst_cellmath__60_0_I279 (.Y(N2856), .A(N2773), .B(N11706));
NOR2XL inst_cellmath__60_0_I280 (.Y(N2673), .A(N2773), .B(N11708));
NOR2XL inst_cellmath__60_0_I281 (.Y(N2820), .A(N2773), .B(N11719));
NOR2XL inst_cellmath__60_0_I282 (.Y(N2635), .A(N2773), .B(N11728));
NOR2XL inst_cellmath__60_0_I283 (.Y(N2776), .A(N2773), .B(N2705));
NOR2XL inst_cellmath__60_0_I284 (.Y(N2593), .A(N2773), .B(N2777));
OR2XL inst_cellmath__60_0_I285 (.Y(N2829), .A(N2773), .B(N2848));
INVXL inst_cellmath__60_0_I286 (.Y(N2609), .A(N11688));
NOR2XL inst_cellmath__60_0_I287 (.Y(N2892), .A(N11688), .B(N11697));
NOR2XL inst_cellmath__60_0_I288 (.Y(N2709), .A(N11688), .B(N11706));
NOR2XL inst_cellmath__60_0_I289 (.Y(N2851), .A(N11688), .B(N11708));
NOR2XL inst_cellmath__60_0_I290 (.Y(N2666), .A(N11688), .B(N11719));
NOR2XL inst_cellmath__60_0_I291 (.Y(N2812), .A(N11688), .B(N11728));
NOR2XL inst_cellmath__60_0_I292 (.Y(N2624), .A(N11688), .B(N2705));
NOR2XL inst_cellmath__60_0_I293 (.Y(N2768), .A(N11688), .B(N2777));
OR2XL inst_cellmath__60_0_I294 (.Y(N2894), .A(N11688), .B(N2848));
INVXL inst_cellmath__60_0_I295 (.Y(N2788), .A(N11697));
NOR2XL inst_cellmath__60_0_I296 (.Y(N2742), .A(N11697), .B(N11706));
NOR2XL inst_cellmath__60_0_I297 (.Y(N2885), .A(N11697), .B(N11708));
NOR2XL inst_cellmath__60_0_I298 (.Y(N2701), .A(N11697), .B(N11719));
NOR2XL inst_cellmath__60_0_I299 (.Y(N2845), .A(N11697), .B(N11728));
NOR2XL inst_cellmath__60_0_I300 (.Y(N2659), .A(N11697), .B(N2705));
NOR2XL inst_cellmath__60_0_I301 (.Y(N2804), .A(N11697), .B(N2777));
OR2XL inst_cellmath__60_0_I302 (.Y(N2642), .A(N11697), .B(N2848));
INVXL inst_cellmath__60_0_I303 (.Y(N2825), .A(N11706));
NOR2XL inst_cellmath__60_0_I304 (.Y(N2780), .A(N11706), .B(N11708));
NOR2XL inst_cellmath__60_0_I305 (.Y(N2597), .A(N11706), .B(N11719));
NOR2XL inst_cellmath__60_0_I306 (.Y(N2735), .A(N11706), .B(N11728));
NOR2XL inst_cellmath__60_0_I307 (.Y(N2879), .A(N11706), .B(N2705));
NOR2XL inst_cellmath__60_0_I308 (.Y(N2694), .A(N11706), .B(N2777));
OR2XL inst_cellmath__60_0_I309 (.Y(N2711), .A(N11706), .B(N2848));
INVXL inst_cellmath__60_0_I310 (.Y(N2712), .A(N11708));
NOR2XL inst_cellmath__60_0_I311 (.Y(N2670), .A(N11708), .B(N11719));
NOR2XL inst_cellmath__60_0_I312 (.Y(N2816), .A(N11708), .B(N11728));
NOR2XL inst_cellmath__60_0_I313 (.Y(N2630), .A(N11708), .B(N2705));
NOR2XL inst_cellmath__60_0_I314 (.Y(N2772), .A(N11708), .B(N2777));
OR2XL inst_cellmath__60_0_I315 (.Y(N2784), .A(N11708), .B(N2848));
INVXL inst_cellmath__60_0_I316 (.Y(N2791), .A(N11719));
NOR2XL inst_cellmath__60_0_I317 (.Y(N2746), .A(N11719), .B(N11728));
NOR2XL inst_cellmath__60_0_I318 (.Y(N2887), .A(N11719), .B(N2705));
NOR2XL inst_cellmath__60_0_I319 (.Y(N2704), .A(N11719), .B(N2777));
OR2XL inst_cellmath__60_0_I320 (.Y(N2853), .A(N11719), .B(N2848));
INVXL inst_cellmath__60_0_I321 (.Y(N2722), .A(N11728));
NOR2XL inst_cellmath__60_0_I322 (.Y(N2681), .A(N11728), .B(N2705));
NOR2XL inst_cellmath__60_0_I323 (.Y(N2831), .A(N11728), .B(N2777));
OR2XL inst_cellmath__60_0_I324 (.Y(N2600), .A(N11728), .B(N2848));
INVXL inst_cellmath__60_0_I325 (.Y(N2843), .A(N2705));
NOR2XL inst_cellmath__60_0_I326 (.Y(N2801), .A(N2705), .B(N2777));
OR2XL inst_cellmath__60_0_I327 (.Y(N2668), .A(N2705), .B(N2848));
INVXL inst_cellmath__60_0_I328 (.Y(N2821), .A(N2777));
ADDHX1 inst_cellmath__60_0_I329 (.CO(N2814), .S(N2739), .A(N11662), .B(N2675));
ADDHX1 inst_cellmath__60_0_I330 (.CO(N2626), .S(N2882), .A(N2629), .B(N2822));
ADDHX1 inst_cellmath__60_0_I331 (.CO(N2770), .S(N2697), .A(N2616), .B(N2636));
ADDFX1 inst_cellmath__60_0_I332 (.CO(N2589), .S(N2842), .A(N2771), .B(N2763), .CI(N2626));
ADDHX1 inst_cellmath__60_0_I333 (.CO(N2726), .S(N2656), .A(N2585), .B(N2779));
ADDFX1 inst_cellmath__60_0_I334 (.CO(N2866), .S(N2800), .A(N2770), .B(N2590), .CI(N2656));
ADDHX1 inst_cellmath__60_0_I335 (.CO(N2684), .S(N2615), .A(N2609), .B(N2595));
ADDFX1 inst_cellmath__60_0_I336 (.CO(N2833), .S(N2755), .A(N2727), .B(N2578), .CI(N2721));
ADDFX1 inst_cellmath__60_0_I337 (.CO(N2645), .S(N2577), .A(N2615), .B(N2726), .CI(N2755));
ADDHX1 inst_cellmath__60_0_I338 (.CO(N2789), .S(N2714), .A(N2715), .B(N2732));
ADDFX1 inst_cellmath__60_0_I339 (.CO(N2605), .S(N2855), .A(N2868), .B(N2862), .CI(N2684));
ADDFX1 inst_cellmath__60_0_I340 (.CO(N2743), .S(N2672), .A(N2833), .B(N2714), .CI(N2855));
ADDHX1 inst_cellmath__60_0_I341 (.CO(N2886), .S(N2819), .A(N2788), .B(N2878));
ADDFX1 inst_cellmath__60_0_I342 (.CO(N2702), .S(N2633), .A(N2685), .B(N2892), .CI(N2680));
ADDFX1 inst_cellmath__60_0_I343 (.CO(N2846), .S(N2775), .A(N2789), .B(N2856), .CI(N2819));
ADDFX1 inst_cellmath__60_0_I344 (.CO(N2660), .S(N2592), .A(N2633), .B(N2605), .CI(N2775));
ADDHX1 inst_cellmath__60_0_I345 (.CO(N2806), .S(N2730), .A(N2709), .B(N2691));
ADDFX1 inst_cellmath__60_0_I346 (.CO(N2619), .S(N2872), .A(N2834), .B(N2673), .CI(N2830));
ADDFX1 inst_cellmath__60_0_I347 (.CO(N2760), .S(N2688), .A(N2730), .B(N2886), .CI(N2702));
ADDFX1 inst_cellmath__60_0_I348 (.CO(N2583), .S(N2837), .A(N2846), .B(N2872), .CI(N2688));
ADDHX1 inst_cellmath__60_0_I349 (.CO(N2719), .S(N2650), .A(N2825), .B(N2839));
ADDFX1 inst_cellmath__60_0_I350 (.CO(N2859), .S(N2794), .A(N2643), .B(N2742), .CI(N2647));
ADDFX1 inst_cellmath__60_0_I351 (.CO(N2677), .S(N2608), .A(N2820), .B(N2851), .CI(N2806));
ADDFX1 inst_cellmath__60_0_I352 (.CO(N2827), .S(N2750), .A(N2650), .B(N2619), .CI(N2794));
ADDFX1 inst_cellmath__60_0_I353 (.CO(N2639), .S(N2891), .A(N2608), .B(N2760), .CI(N2750));
XNOR2X1 inst_cellmath__60_0_I354 (.Y(N2708), .A(N2885), .B(N2790));
OR2XL inst_cellmath__60_0_I355 (.Y(N2782), .A(N2885), .B(N2790));
ADDFX1 inst_cellmath__60_0_I356 (.CO(N2736), .S(N2665), .A(N2785), .B(N2666), .CI(N2635));
ADDFX1 inst_cellmath__60_0_I357 (.CO(N2880), .S(N2810), .A(N2719), .B(N2611), .CI(N2708));
ADDFX1 inst_cellmath__60_0_I358 (.CO(N2695), .S(N2623), .A(N2677), .B(N2859), .CI(N2665));
ADDFX1 inst_cellmath__60_0_I359 (.CO(N2841), .S(N2767), .A(N2827), .B(N2810), .CI(N2623));
ADDFX1 inst_cellmath__60_0_I360 (.CO(N2655), .S(N2587), .A(N2780), .B(N2712), .CI(N2602));
ADDFX1 inst_cellmath__60_0_I361 (.CO(N2798), .S(N2724), .A(N2776), .B(N2701), .CI(N2812));
ADDFX1 inst_cellmath__60_0_I362 (.CO(N2614), .S(N2865), .A(N2782), .B(N2679), .CI(N2736));
ADDFX1 inst_cellmath__60_0_I363 (.CO(N2754), .S(N2683), .A(N2724), .B(N2587), .CI(N2880));
ADDFX1 inst_cellmath__60_0_I364 (.CO(N2896), .S(N2832), .A(N2695), .B(N2865), .CI(N2683));
ADDFX1 inst_cellmath__60_0_I365 (.CO(N2713), .S(N2644), .A(N2593), .B(N2597), .CI(N2624));
ADDFX1 inst_cellmath__60_0_I366 (.CO(N2854), .S(N2787), .A(N2753), .B(N2845), .CI(N2655));
ADDFX1 inst_cellmath__60_0_I367 (.CO(N2671), .S(N2604), .A(N2644), .B(N2798), .CI(N2614));
ADDFX1 inst_cellmath__60_0_I368 (.CO(N2817), .S(N2741), .A(N2754), .B(N2787), .CI(N2604));
ADDFX1 inst_cellmath__60_0_I369 (.CO(N2632), .S(N2884), .A(N2670), .B(N2791), .CI(N2768));
ADDFX1 inst_cellmath__60_0_I370 (.CO(N2774), .S(N2699), .A(N2659), .B(N2735), .CI(N2829));
ADDFX1 inst_cellmath__60_0_I371 (.CO(N2591), .S(N2844), .A(N2884), .B(N2713), .CI(N2699));
ADDFX1 inst_cellmath__60_0_I372 (.CO(N2729), .S(N2658), .A(N2671), .B(N2854), .CI(N2844));
ADDFX1 inst_cellmath__60_0_I373 (.CO(N2870), .S(N2802), .A(N2804), .B(N2816), .CI(N2879));
ADDFX1 inst_cellmath__60_0_I374 (.CO(N2686), .S(N2617), .A(N2632), .B(N2894), .CI(N2774));
ADDFX1 inst_cellmath__60_0_I375 (.CO(N2835), .S(N2758), .A(N2591), .B(N2802), .CI(N2617));
ADDFX1 inst_cellmath__60_0_I376 (.CO(N2649), .S(N2581), .A(N2746), .B(N2722), .CI(N2694));
ADDFX1 inst_cellmath__60_0_I377 (.CO(N2792), .S(N2717), .A(N2642), .B(N2630), .CI(N2870));
ADDFX1 inst_cellmath__60_0_I378 (.CO(N2606), .S(N2858), .A(N2686), .B(N2581), .CI(N2717));
ADDFX1 inst_cellmath__60_0_I379 (.CO(N2748), .S(N2674), .A(N2772), .B(N2887), .CI(N2711));
ADDFX1 inst_cellmath__60_0_I380 (.CO(N2889), .S(N2824), .A(N2674), .B(N2649), .CI(N2792));
ADDFX1 inst_cellmath__60_0_I381 (.CO(N2706), .S(N2638), .A(N2681), .B(N2843), .CI(N2704));
ADDFX1 inst_cellmath__60_0_I382 (.CO(N2849), .S(N2778), .A(N2748), .B(N2784), .CI(N2638));
ADDFX1 inst_cellmath__60_0_I383 (.CO(N2663), .S(N2596), .A(N2853), .B(N2831), .CI(N2706));
ADDFX1 inst_cellmath__60_0_I384 (.CO(N2809), .S(N2734), .A(N2801), .B(N2821), .CI(N2600));
AND2XL inst_cellmath__60_0_I387 (.Y(N2764), .A(N2815), .B(N2739));
NAND2XL inst_cellmath__60_0_I389 (.Y(N2586), .A(N2814), .B(N2882));
AND2XL inst_cellmath__60_0_I391 (.Y(N2723), .A(N2697), .B(N2842));
NOR2XL inst_cellmath__60_0_I392 (.Y(N2797), .A(N2589), .B(N2800));
NAND2XL inst_cellmath__60_0_I393 (.Y(N2863), .A(N2589), .B(N2800));
AND2XL inst_cellmath__60_0_I395 (.Y(N2682), .A(N2866), .B(N2577));
NOR4X1 inst_cellmath__60_0_I5075 (.Y(N2895), .A(N2876), .B(N11661), .C(N11660), .D(N11670));
OAI22XL inst_cellmath__60_0_I5047 (.Y(N2628), .A0(N2764), .A1(N2895), .B0(N2815), .B1(N2739));
AOI2BB2X1 inst_cellmath__60_0_I5048 (.Y(N2869), .A0N(N2814), .A1N(N2882), .B0(N2628), .B1(N2586));
OAI22XL inst_cellmath__60_0_I5049 (.Y(N2745), .A0(N2723), .A1(N2869), .B0(N2697), .B1(N2842));
AOI21XL inst_cellmath__60_0_I404 (.Y(N2621), .A0(N2863), .A1(N2745), .B0(N2797));
OAI22XL inst_cellmath__60_0_I5050 (.Y(N2847), .A0(N2682), .A1(N2621), .B0(N2866), .B1(N2577));
NOR2XL inst_cellmath__60_0_I420 (.Y(N2661), .A(N2645), .B(N2672));
XOR2XL inst_cellmath__60_0_I421 (.Y(N2731), .A(N2645), .B(N2672));
XOR2XL inst_cellmath__60_0_I423 (.Y(N2875), .A(N2743), .B(N2592));
XOR2XL inst_cellmath__60_0_I425 (.Y(N2689), .A(N2660), .B(N2837));
NOR2XL inst_cellmath__60_0_I426 (.Y(N2762), .A(N2583), .B(N2891));
XOR2XL inst_cellmath__60_0_I427 (.Y(N2838), .A(N2583), .B(N2891));
NOR2XL inst_cellmath__60_0_I428 (.Y(N2584), .A(N2639), .B(N2767));
XOR2XL inst_cellmath__60_0_I429 (.Y(N2652), .A(N2639), .B(N2767));
NOR2XL inst_cellmath__60_0_I430 (.Y(N2720), .A(N2841), .B(N2832));
XOR2XL inst_cellmath__60_0_I431 (.Y(N2795), .A(N2841), .B(N2832));
NOR2XL inst_cellmath__60_0_I432 (.Y(N2861), .A(N2896), .B(N2741));
XOR2XL inst_cellmath__60_0_I433 (.Y(N2610), .A(N2896), .B(N2741));
NOR2XL inst_cellmath__60_0_I434 (.Y(N2678), .A(N2817), .B(N2658));
XOR2XL inst_cellmath__60_0_I435 (.Y(N2752), .A(N2817), .B(N2658));
NOR2XL inst_cellmath__60_0_I436 (.Y(N2828), .A(N2729), .B(N2758));
XOR2XL inst_cellmath__60_0_I437 (.Y(N2893), .A(N2729), .B(N2758));
NOR2XL inst_cellmath__60_0_I438 (.Y(N2641), .A(N2835), .B(N2858));
XOR2XL inst_cellmath__60_0_I439 (.Y(N2710), .A(N2835), .B(N2858));
NOR2XL inst_cellmath__60_0_I440 (.Y(N2783), .A(N2824), .B(N2606));
XOR2XL inst_cellmath__60_0_I441 (.Y(N2852), .A(N2824), .B(N2606));
NOR2XL inst_cellmath__60_0_I442 (.Y(N2599), .A(N2889), .B(N2778));
XOR2XL inst_cellmath__60_0_I443 (.Y(N2667), .A(N2889), .B(N2778));
NOR2XL inst_cellmath__60_0_I444 (.Y(N2738), .A(N2596), .B(N2849));
XOR2XL inst_cellmath__60_0_I445 (.Y(N2813), .A(N2596), .B(N2849));
NOR2XL inst_cellmath__60_0_I446 (.Y(N2881), .A(N2734), .B(N2663));
XOR2XL inst_cellmath__60_0_I447 (.Y(N2625), .A(N2734), .B(N2663));
NOR2XL inst_cellmath__60_0_I448 (.Y(N2696), .A(N2668), .B(N2809));
XOR2XL inst_cellmath__60_0_I449 (.Y(N2769), .A(N2668), .B(N2809));
NAND2BXL inst_cellmath__60_0_I450 (.Y(N2588), .AN(N2848), .B(N2777));
AO21XL inst_cellmath__60_0_I451 (.Y(N2799), .A0(N2731), .A1(N2847), .B0(N2661));
OR2XL gen2_alt_A_I14169 (.Y(N11749), .A(N2743), .B(N2592));
OAI2BB1X1 gen2_alt_A_I5092 (.Y(N2576), .A0N(N2875), .A1N(N2799), .B0(N11749));
OR2XL gena_A_I14170 (.Y(N11756), .A(N2660), .B(N2837));
NAND2XL gena_A_I5094 (.Y(N11758), .A(N2689), .B(N2576));
NAND2XL gena_A_I5095 (.Y(N2818), .A(N11756), .B(N11758));
AO21XL inst_cellmath__60_0_I454 (.Y(N2871), .A0(N2838), .A1(N2818), .B0(N2762));
AO21XL inst_cellmath__60_0_I455 (.Y(N2749), .A0(N2652), .A1(N2871), .B0(N2584));
AO21XL inst_cellmath__60_0_I456 (.Y(N2766), .A0(N2795), .A1(N2749), .B0(N2720));
AO21XL inst_cellmath__60_0_I457 (.Y(N2603), .A0(N2610), .A1(N2766), .B0(N2861));
AO21XL inst_cellmath__60_0_I458 (.Y(N2580), .A0(N2752), .A1(N2603), .B0(N2678));
AO21XL inst_cellmath__60_0_I459 (.Y(N2690), .A0(N2893), .A1(N2580), .B0(N2828));
AO21XL inst_cellmath__60_0_I460 (.Y(N2627), .A0(N2710), .A1(N2690), .B0(N2641));
AO21XL inst_cellmath__60_0_I461 (.Y(N2703), .A0(N2852), .A1(N2627), .B0(N2783));
AO21XL inst_cellmath__60_0_I462 (.Y(N2601), .A0(N2667), .A1(N2703), .B0(N2599));
AO21XL inst_cellmath__60_0_I463 (.Y(N2634), .A0(N2813), .A1(N2601), .B0(N2738));
AO21XL inst_cellmath__60_0_I464 (.Y(N2811), .A0(N2625), .A1(N2634), .B0(N2881));
AO21XL inst_cellmath__60_0_I465 (.Y(N2803), .A0(N2769), .A1(N2811), .B0(N2696));
XNOR2X1 inst_cellmath__60_0_I478 (.Y(inst_cellmath__60[21]), .A(N2601), .B(N2813));
XNOR2X1 inst_cellmath__60_0_I479 (.Y(inst_cellmath__60[22]), .A(N2634), .B(N2625));
CLKXOR2X1 inst_cellmath__60_0_I480 (.Y(inst_cellmath__60[23]), .A(N2811), .B(N2769));
XNOR2X1 inst_cellmath__60_0_I481 (.Y(inst_cellmath__60[24]), .A(N2803), .B(N2588));
INVXL cynw_cm_float_rcp_I482 (.Y(N3346), .A(a_man[16]));
INVXL cynw_cm_float_rcp_I483 (.Y(N3723), .A(a_man[17]));
AOI22X1 cynw_cm_float_rcp_I484 (.Y(N3482), .A0(N3346), .A1(a_man[17]), .B0(N3723), .B1(a_man[16]));
NAND2X1 cynw_cm_float_rcp_I485 (.Y(N3869), .A(N3723), .B(N3346));
NAND2X1 cynw_cm_float_rcp_I486 (.Y(N3344), .A(N3723), .B(a_man[16]));
NOR2X1 cynw_cm_float_rcp_I487 (.Y(N3752), .A(N3723), .B(N3346));
NAND2X1 cynw_cm_float_rcp_I488 (.Y(N3222), .A(a_man[16]), .B(a_man[17]));
NOR2X1 cynw_cm_float_rcp_I489 (.Y(N3636), .A(N3723), .B(a_man[16]));
NOR2XL cynw_cm_float_rcp_I490 (.Y(N4036), .A(a_man[17]), .B(a_man[16]));
NOR2X1 cynw_cm_float_rcp_I491 (.Y(N3517), .A(a_man[17]), .B(N3346));
INVX2 cynw_cm_float_rcp_I492 (.Y(N3641), .A(a_man[18]));
AOI22XL cynw_cm_float_rcp_I493 (.Y(N3923), .A0(N3641), .A1(N3869), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I494 (.Y(N3857), .A0(N3641), .A1(N3636), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I495 (.Y(N4058), .A0(N3641), .A1(N3222), .B0(N3869), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I496 (.Y(N3390), .A(a_man[18]), .B(N3752));
AOI22XL cynw_cm_float_rcp_I497 (.Y(N3382), .A0(N3641), .A1(N3752), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I498 (.Y(N3583), .A0(N3641), .A1(N3723), .B0(a_man[16]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I499 (.Y(N3789), .A(N3344));
AOI22XL cynw_cm_float_rcp_I500 (.Y(N3802), .A0(N3641), .A1(N3344), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I501 (.Y(N3269), .A0(N3641), .A1(a_man[17]), .B0(a_man[16]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I502 (.Y(N3488), .A(N3482));
AOI22XL cynw_cm_float_rcp_I503 (.Y(N3672), .A0(N3641), .A1(N3636), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I504 (.Y(N4091), .A0(N3641), .A1(N3723), .B0(N3752), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I505 (.Y(N4073), .A(N3641), .B(N3222));
AOI22XL cynw_cm_float_rcp_I506 (.Y(N3600), .A0(N3641), .A1(N3636), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I507 (.Y(N4003), .A0(N3641), .A1(a_man[16]), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I508 (.Y(N3562), .A0(N3641), .A1(N3222), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I509 (.Y(N3969), .A0(N3641), .A1(N4036), .B0(a_man[17]), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I510 (.Y(N3689), .A(a_man[18]), .B(N3636));
AOI22XL cynw_cm_float_rcp_I511 (.Y(N3364), .A0(N3641), .A1(a_man[16]), .B0(N3869), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I512 (.Y(N3565), .A(N3641), .B(N3752));
NOR2XL cynw_cm_float_rcp_I513 (.Y(N3442), .A(a_man[18]), .B(N3517));
AOI22XL cynw_cm_float_rcp_I515 (.Y(N3535), .A0(N3641), .A1(N3723), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I516 (.Y(N3736), .A0(N3641), .A1(N3752), .B0(N3869), .B1(a_man[18]));
NAND2X1 cynw_cm_float_rcp_I517 (.Y(N3708), .A(N3346), .B(a_man[17]));
AOI22X1 cynw_cm_float_rcp_I518 (.Y(N3465), .A0(a_man[16]), .A1(a_man[17]), .B0(N3723), .B1(N3346));
NOR2XL cynw_cm_float_rcp_I519 (.Y(N4137), .A(N3641), .B(N4036));
AOI22XL cynw_cm_float_rcp_I520 (.Y(N3614), .A0(N3641), .A1(a_man[17]), .B0(N3723), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I521 (.Y(N4015), .A(a_man[17]), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I522 (.Y(N3494), .A0(N3641), .A1(N3465), .B0(N3708), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I523 (.Y(N3486), .A(N3641), .B(N3346));
AOI22XL cynw_cm_float_rcp_I524 (.Y(N3891), .A0(N3641), .A1(N3482), .B0(N3222), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I525 (.Y(N4099), .A0(N3641), .A1(N3222), .B0(N3465), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I526 (.Y(N3369), .A0(N3641), .A1(N3752), .B0(N3465), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I527 (.Y(N3899), .A0(N3641), .A1(a_man[16]), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I528 (.Y(N3244), .A0(N3641), .A1(N3465), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I529 (.Y(N3450), .A0(N3641), .A1(N3708), .B0(N3517), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I530 (.Y(N3395), .A(N3465));
AOI22XL cynw_cm_float_rcp_I531 (.Y(N3779), .A0(N3641), .A1(N3869), .B0(N4036), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I532 (.Y(N3250), .A(a_man[18]), .B(N3869));
NAND2XL cynw_cm_float_rcp_I533 (.Y(N3666), .A(N3641), .B(N4036));
NAND2XL cynw_cm_float_rcp_I534 (.Y(N3910), .A(N3346), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I535 (.Y(N4065), .A0(N3641), .A1(a_man[17]), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I536 (.Y(N3585), .A0(N3641), .A1(N4036), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I537 (.Y(N3543), .A0(N3641), .A1(a_man[17]), .B0(N3517), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I538 (.Y(N3989), .A(N3641), .B(a_man[17]));
NAND2XL cynw_cm_float_rcp_I539 (.Y(N3463), .A(N3641), .B(a_man[16]));
AOI22XL cynw_cm_float_rcp_I540 (.Y(N3347), .A0(N3641), .A1(N3869), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I541 (.Y(N3548), .A0(N3641), .A1(a_man[17]), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I542 (.Y(N3754), .A0(N3641), .A1(N3636), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I543 (.Y(N3949), .A0(N3641), .A1(a_man[17]), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I544 (.Y(N3429), .A0(N3641), .A1(N3465), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I545 (.Y(N3638), .A0(N3641), .A1(N3752), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I546 (.Y(N3419), .A0(N3641), .A1(N3346), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I547 (.Y(N3830), .A0(N3641), .A1(N3482), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I548 (.Y(N3301), .A0(N3641), .A1(N4036), .B0(N3869), .B1(a_man[18]));
CLKINVX6 cynw_cm_float_rcp_I551 (.Y(N3714), .A(a_man[19]));
AOI22XL cynw_cm_float_rcp_I552 (.Y(N3770), .A0(N3714), .A1(N4137), .B0(N3923), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I553 (.Y(N3971), .A0(N3714), .A1(N3346), .B0(N3857), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I555 (.Y(N3240), .A0(N3714), .A1(a_man[17]), .B0(N4058), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I556 (.Y(N3447), .A0(N3714), .A1(N3614), .B0(N3390), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I557 (.Y(N3655), .A(N3714), .B(N4015));
AOI22XL cynw_cm_float_rcp_I558 (.Y(N3407), .A0(N3714), .A1(N3494), .B0(N3382), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I559 (.Y(N3619), .A0(N3714), .A1(N3486), .B0(N3583), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I560 (.Y(N3821), .A0(N3714), .A1(N3891), .B0(N3789), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I561 (.Y(N4020), .A0(N3714), .A1(N4099), .B0(N3802), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I562 (.Y(N3291), .A0(N3714), .A1(N3369), .B0(N3269), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I563 (.Y(N3500), .A0(N3714), .A1(N3899), .B0(N3488), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I564 (.Y(N3704), .A0(N3714), .A1(N3269), .B0(N3672), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I565 (.Y(N3906), .A0(N3714), .A1(N3899), .B0(N4091), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I566 (.Y(N4113), .A0(N3714), .A1(N3244), .B0(N4073), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I567 (.Y(N3380), .A0(N3714), .A1(N3450), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I568 (.Y(N3579), .A0(N3714), .A1(N3395), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I569 (.Y(N3783), .A0(N3714), .A1(N3779), .B0(a_man[18]), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I570 (.Y(N3984), .A(a_man[19]), .B(N3250));
NOR2XL cynw_cm_float_rcp_I571 (.Y(N3711), .A(a_man[19]), .B(N3666));
AOI22XL cynw_cm_float_rcp_I572 (.Y(N3836), .A0(N3714), .A1(N2381), .B0(N3600), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I573 (.Y(N4034), .A0(N3714), .A1(N3910), .B0(N3802), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I574 (.Y(N3308), .A0(N3714), .A1(N4065), .B0(N4003), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I575 (.Y(N3515), .A0(N3714), .A1(N3585), .B0(N3562), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I576 (.Y(N3718), .A0(N3714), .A1(N3543), .B0(N3969), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I577 (.Y(N3922), .A0(N3714), .A1(N3989), .B0(N3689), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I578 (.Y(N4124), .A0(N3714), .A1(N3463), .B0(N3364), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I579 (.Y(N3388), .A0(N3714), .A1(N3969), .B0(N3565), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I580 (.Y(N3594), .A0(N3714), .A1(N4065), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I581 (.Y(N3800), .A0(N3714), .A1(N3347), .B0(N2381), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I582 (.Y(N3997), .A0(N3714), .A1(N3548), .B0(N3488), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I583 (.Y(N3267), .A0(N3714), .A1(N3754), .B0(N3535), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I584 (.Y(N3476), .A0(N3714), .A1(N3543), .B0(N3736), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I585 (.Y(N3684), .A0(N3714), .A1(N3949), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I586 (.Y(N3883), .A0(N3714), .A1(N3429), .B0(N2381), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I587 (.Y(N4089), .A(N3714), .B(N3638));
NOR2XL cynw_cm_float_rcp_I588 (.Y(N3560), .A(a_man[19]), .B(N4137));
AOI22XL cynw_cm_float_rcp_I589 (.Y(N3236), .A0(N3714), .A1(N3419), .B0(N3346), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I590 (.Y(N3441), .A0(N3714), .A1(N3830), .B0(N3723), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I591 (.Y(N3650), .A0(N3714), .A1(N3301), .B0(N3641), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I592 (.Y(N3850), .A(N3714), .B(N3666));
NAND2XL cynw_cm_float_rcp_I593 (.Y(N3326), .A(N3714), .B(N3250));
NOR2XL cynw_cm_float_rcp_I594 (.Y(N4120), .A(N3641), .B(N3723));
AOI22XL cynw_cm_float_rcp_I595 (.Y(N3590), .A0(N3641), .A1(N3869), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I596 (.Y(N3992), .A0(N3641), .A1(N3636), .B0(N3517), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I597 (.Y(N3757), .A0(N3641), .A1(N3222), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I598 (.Y(N3957), .A0(N3641), .A1(N4036), .B0(a_man[16]), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I599 (.Y(N4041), .A(a_man[18]), .B(N4036));
AOI22XL cynw_cm_float_rcp_I600 (.Y(N3469), .A0(N3641), .A1(a_man[16]), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I601 (.Y(N3876), .A0(N3641), .A1(N3465), .B0(N3723), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I602 (.Y(N3352), .A0(N3641), .A1(N3708), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I603 (.Y(N3761), .A0(N3641), .A1(N3482), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I604 (.Y(N3229), .A0(N3641), .A1(N3752), .B0(N3723), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I605 (.Y(N3643), .A(N3641), .B(N3222));
AOI22XL cynw_cm_float_rcp_I606 (.Y(N3773), .A0(N3641), .A1(a_man[16]), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I607 (.Y(N3973), .A0(N3641), .A1(N3517), .B0(N3222), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I608 (.Y(N3242), .A(N3641), .B(N3869));
NOR2XL cynw_cm_float_rcp_I609 (.Y(N3856), .A(a_man[18]), .B(N3222));
AOI22XL cynw_cm_float_rcp_I610 (.Y(N4046), .A0(N3641), .A1(N3465), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I611 (.Y(N3940), .A0(N3641), .A1(N3708), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I612 (.Y(N3526), .A0(N3641), .A1(N3344), .B0(N3465), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I613 (.Y(N3705), .A0(N3641), .A1(N3708), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I614 (.Y(N3933), .A0(N3641), .A1(N3752), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I615 (.Y(N3399), .A0(N3641), .A1(N3517), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I616 (.Y(N3811), .A0(N3641), .A1(a_man[16]), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I617 (.Y(N3787), .A0(N3641), .A1(N3723), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I618 (.Y(N3279), .A0(N3641), .A1(N3723), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I619 (.Y(N3351), .A0(N3641), .A1(N3346), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I620 (.Y(N4134), .A0(N3641), .A1(N3752), .B0(N3222), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I621 (.Y(N3693), .A0(N3641), .A1(N3869), .B0(N3723), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I622 (.Y(N3608), .A(N3869));
AOI22XL cynw_cm_float_rcp_I623 (.Y(N3810), .A0(N3641), .A1(N3517), .B0(N3752), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I624 (.Y(N4008), .A(N4036), .B(a_man[18]));
NAND2XL cynw_cm_float_rcp_I625 (.Y(N4102), .A(N3641), .B(N3708));
AOI22XL cynw_cm_float_rcp_I626 (.Y(N3893), .A0(N3641), .A1(N3723), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I627 (.Y(N4101), .A0(N3641), .A1(N3723), .B0(N3465), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I628 (.Y(N3570), .A0(N3641), .A1(N3636), .B0(N3465), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I629 (.Y(N3976), .A0(N3641), .A1(N3344), .B0(N3517), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I630 (.Y(N3452), .A(N3869), .B(a_man[18]));
NOR2XL cynw_cm_float_rcp_I631 (.Y(N3624), .A(N3641), .B(a_man[16]));
NAND2XL cynw_cm_float_rcp_I632 (.Y(N3505), .A(N3641), .B(N3344));
AOI22XL cynw_cm_float_rcp_I633 (.Y(N3587), .A0(N3641), .A1(a_man[16]), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I634 (.Y(N3794), .A0(N3641), .A1(N3752), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I635 (.Y(N3466), .A0(N3641), .A1(N3708), .B0(N3222), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I636 (.Y(N3874), .A(N3641), .B(N3517));
AOI22XL cynw_cm_float_rcp_I637 (.Y(N3860), .A0(N3641), .A1(N3708), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I638 (.Y(N3929), .A0(N3641), .A1(a_man[17]), .B0(N3465), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I639 (.Y(N3335), .A(N3641), .B(N3752));
NAND2XL cynw_cm_float_rcp_I640 (.Y(N3243), .A(N3714), .B(N3989));
AOI22XL cynw_cm_float_rcp_I641 (.Y(N3658), .A0(N3714), .A1(N3351), .B0(N3346), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I642 (.Y(N3858), .A0(N3714), .A1(N3876), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I643 (.Y(N4059), .A0(N3714), .A1(N3229), .B0(N3614), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I644 (.Y(N3333), .A0(N3714), .A1(N4015), .B0(N4120), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I645 (.Y(N3538), .A(N3714), .B(N4015));
AOI22XL cynw_cm_float_rcp_I646 (.Y(N3294), .A0(N3714), .A1(N4134), .B0(N3590), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I647 (.Y(N3503), .A0(N3714), .A1(N3693), .B0(N3992), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I648 (.Y(N3707), .A0(N3714), .A1(N3608), .B0(N3757), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I649 (.Y(N3909), .A0(N3714), .A1(N3810), .B0(N3957), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I650 (.Y(N4116), .A0(N3714), .A1(N4008), .B0(N3562), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I651 (.Y(N3383), .A0(N3714), .A1(N4102), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I652 (.Y(N3584), .A0(N3714), .A1(N3893), .B0(N4041), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I653 (.Y(N3790), .A0(N3714), .A1(N4101), .B0(N3469), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I654 (.Y(N3988), .A0(N3714), .A1(N3429), .B0(N3876), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I655 (.Y(N3258), .A0(N3714), .A1(N3570), .B0(N3352), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I656 (.Y(N3462), .A0(N3714), .A1(N3976), .B0(N3761), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I657 (.Y(N3673), .A0(N3714), .A1(N3279), .B0(N3229), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I658 (.Y(N3872), .A0(N3714), .A1(N3452), .B0(N3643), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I659 (.Y(N3743), .A(N3714), .B(N3452));
AOI22XL cynw_cm_float_rcp_I660 (.Y(N3314), .A0(N3714), .A1(N3624), .B0(N3773), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I661 (.Y(N3521), .A0(N3714), .A1(N4046), .B0(N3973), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I662 (.Y(N3722), .A0(N3714), .A1(N3505), .B0(N3242), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I663 (.Y(N3927), .A0(N3714), .A1(N4137), .B0(N3856), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I664 (.Y(N4130), .A0(N3714), .A1(N3587), .B0(N3802), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I665 (.Y(N3393), .A0(N3714), .A1(N3794), .B0(N4046), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I666 (.Y(N3602), .A0(N3714), .A1(N3347), .B0(N3940), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I667 (.Y(N3807), .A0(N3714), .A1(N3590), .B0(N3562), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I668 (.Y(N4004), .A0(N3714), .A1(N3466), .B0(N4091), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I669 (.Y(N3274), .A0(N3714), .A1(N3811), .B0(N3526), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I670 (.Y(N3481), .A0(N3714), .A1(N3874), .B0(N3526), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I671 (.Y(N3690), .A(N3714), .B(N3860));
AOI22XL cynw_cm_float_rcp_I672 (.Y(N4095), .A0(N3714), .A1(N3923), .B0(N3957), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I673 (.Y(N3365), .A0(N3714), .A1(a_man[17]), .B0(N3705), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I674 (.Y(N3566), .A0(N3714), .A1(N2381), .B0(N3933), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I675 (.Y(N3769), .A0(N3714), .A1(N3346), .B0(N3399), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I676 (.Y(N3970), .A0(N3714), .A1(N3723), .B0(N4065), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I677 (.Y(N3238), .A0(N3714), .A1(N3469), .B0(N3811), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I678 (.Y(N3445), .A0(N3714), .A1(N3929), .B0(N3787), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I679 (.Y(N3653), .A0(N3714), .A1(N3335), .B0(N3279), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I680 (.Y(N3854), .A0(N3714), .A1(a_man[18]), .B0(N2381), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I681 (.Y(N4054), .A(a_man[19]), .B(a_man[18]));
NAND2XL cynw_cm_float_rcp_I682 (.Y(N3737), .A(N3714), .B(N3641));
INVX3 cynw_cm_float_rcp_I683 (.Y(N3411), .A(a_man[20]));
AOI22XL cynw_cm_float_rcp_I684 (.Y(N3820), .A0(N3411), .A1(N3243), .B0(N3770), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I685 (.Y(N4019), .A0(N3411), .A1(N3658), .B0(N3971), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I686 (.Y(N3290), .A0(N3411), .A1(N3858), .B0(N3240), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I687 (.Y(N3499), .A0(N3411), .A1(N4059), .B0(N3447), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I688 (.Y(N3702), .A0(N3411), .A1(N3333), .B0(N3655), .B1(a_man[20]));
NOR2XL cynw_cm_float_rcp_I689 (.Y(N3904), .A(a_man[20]), .B(N3538));
AOI22XL cynw_cm_float_rcp_I690 (.Y(N4069), .A0(N3411), .A1(N3294), .B0(N3407), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I691 (.Y(N3341), .A0(N3411), .A1(N3503), .B0(N3619), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I692 (.Y(N3546), .A0(N3411), .A1(N3707), .B0(N3821), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I693 (.Y(N3749), .A0(N3411), .A1(N3909), .B0(N4020), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I694 (.Y(N3952), .A0(N3411), .A1(N4116), .B0(N3291), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I695 (.Y(N3220), .A0(N3411), .A1(N3383), .B0(N3500), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I696 (.Y(N3425), .A0(N3411), .A1(N3584), .B0(N3704), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I697 (.Y(N3634), .A0(N3411), .A1(N3790), .B0(N3906), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I698 (.Y(N3835), .A0(N3411), .A1(N3988), .B0(N4113), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I699 (.Y(N4033), .A0(N3411), .A1(N3258), .B0(N3380), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I700 (.Y(N3306), .A0(N3411), .A1(N3462), .B0(N3579), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I701 (.Y(N3513), .A0(N3411), .A1(N3673), .B0(N3783), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I702 (.Y(N3716), .A0(N3411), .A1(N3872), .B0(N3984), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I703 (.Y(N3920), .A0(N3411), .A1(N3743), .B0(N3711), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I704 (.Y(N4122), .A(N3411), .B(N3560));
AOI22XL cynw_cm_float_rcp_I705 (.Y(N3474), .A0(N3411), .A1(N3314), .B0(N3836), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I706 (.Y(N3682), .A0(N3411), .A1(N3521), .B0(N4034), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I707 (.Y(N3881), .A0(N3411), .A1(N3722), .B0(N3308), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I708 (.Y(N4087), .A0(N3411), .A1(N3927), .B0(N3515), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I709 (.Y(N3357), .A0(N3411), .A1(N4130), .B0(N3718), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I710 (.Y(N3558), .A0(N3411), .A1(N3393), .B0(N3922), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I711 (.Y(N3766), .A0(N3411), .A1(N3602), .B0(N4124), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I712 (.Y(N3967), .A0(N3411), .A1(N3807), .B0(N3388), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I713 (.Y(N3234), .A0(N3411), .A1(N4004), .B0(N3594), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I714 (.Y(N3439), .A0(N3411), .A1(N3274), .B0(N3800), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I715 (.Y(N3648), .A0(N3411), .A1(N3481), .B0(N3997), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I716 (.Y(N3847), .A0(N3411), .A1(N3690), .B0(N3267), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I717 (.Y(N4051), .A0(N3411), .A1(N4095), .B0(N3476), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I718 (.Y(N3325), .A0(N3411), .A1(N3365), .B0(N3684), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I719 (.Y(N3532), .A0(N3411), .A1(N3566), .B0(N3883), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I720 (.Y(N3732), .A0(N3411), .A1(N3769), .B0(N4089), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I721 (.Y(N3936), .A0(N3411), .A1(N3970), .B0(N3560), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I722 (.Y(N4136), .A0(N3411), .A1(N3238), .B0(N3236), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I723 (.Y(N3401), .A0(N3411), .A1(N3445), .B0(N3441), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I724 (.Y(N3612), .A0(N3411), .A1(N3653), .B0(N3650), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I725 (.Y(N3814), .A0(N3411), .A1(N3854), .B0(N3850), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I726 (.Y(N4012), .A0(N3411), .A1(N4054), .B0(N3326), .B1(a_man[20]));
NOR2XL cynw_cm_float_rcp_I727 (.Y(N3283), .A(a_man[20]), .B(N3737));
AOI22XL cynw_cm_float_rcp_I728 (.Y(N3212), .A0(N3641), .A1(N3517), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I729 (.Y(N3792), .A0(N3641), .A1(N3708), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I730 (.Y(N3639), .A0(N3641), .A1(N3752), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I731 (.Y(N3625), .A0(N3641), .A1(N3708), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I732 (.Y(N3315), .A0(N3641), .A1(N3346), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I733 (.Y(N3522), .A0(N3641), .A1(N3752), .B0(N3708), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I734 (.Y(N3724), .A(N3641), .B(N3465));
AOI22XL cynw_cm_float_rcp_I735 (.Y(N3394), .A0(N3641), .A1(N3346), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I736 (.Y(N4025), .A0(N3641), .A1(N3465), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I737 (.Y(N3506), .A0(N3641), .A1(N3344), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I738 (.Y(N3913), .A0(N3641), .A1(a_man[17]), .B0(N3222), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I739 (.Y(N3384), .A(N3641), .B(N3723));
NOR2XL cynw_cm_float_rcp_I740 (.Y(N3739), .A(N3641), .B(N3517));
AOI22XL cynw_cm_float_rcp_I741 (.Y(N4021), .A0(N3641), .A1(N3708), .B0(N3723), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I742 (.Y(N3795), .A0(N3641), .A1(a_man[17]), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I743 (.Y(N3501), .A0(N3641), .A1(N3465), .B0(N3222), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I744 (.Y(N3581), .A0(N3641), .A1(N3708), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I745 (.Y(N3785), .A0(N3641), .A1(a_man[16]), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I746 (.Y(N3985), .A0(N3641), .A1(N3708), .B0(N4036), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I747 (.Y(N3255), .A(N3636));
AOI22XL cynw_cm_float_rcp_I748 (.Y(N3260), .A0(N3641), .A1(a_man[16]), .B0(N3465), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I749 (.Y(N3676), .A0(N3641), .A1(N3482), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I750 (.Y(N3808), .A0(N3641), .A1(N3482), .B0(N3517), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I751 (.Y(N4079), .A0(N3641), .A1(N3482), .B0(N3723), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I752 (.Y(N3489), .A0(N3641), .A1(N3346), .B0(N3636), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I753 (.Y(N3825), .A(N3641), .B(N3465));
NAND2XL cynw_cm_float_rcp_I754 (.Y(N3298), .A(N3708), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I755 (.Y(N3912), .A0(N3641), .A1(N4036), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I756 (.Y(N3586), .A0(N3641), .A1(N4036), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I757 (.Y(N3793), .A0(N3641), .A1(N3465), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I758 (.Y(N3990), .A0(N3641), .A1(N3723), .B0(N3636), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I759 (.Y(N4078), .A(N3222));
NOR2XL cynw_cm_float_rcp_I760 (.Y(N3550), .A(N3641), .B(a_man[17]));
AOI22XL cynw_cm_float_rcp_I761 (.Y(N3958), .A0(N3641), .A1(N3346), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I762 (.Y(N4042), .A0(N3641), .A1(N3723), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I763 (.Y(N3431), .A0(N3641), .A1(a_man[16]), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I764 (.Y(N3889), .A0(N3714), .A1(N3506), .B0(N3212), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I765 (.Y(N4097), .A0(N3714), .A1(N4101), .B0(N3494), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I766 (.Y(N3367), .A0(N3714), .A1(N3811), .B0(N3792), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I767 (.Y(N3568), .A0(N3714), .A1(N3795), .B0(N3279), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I768 (.Y(N3741), .A0(N3714), .A1(N3301), .B0(N3639), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I769 (.Y(N3942), .A0(N3714), .A1(N3736), .B0(N3860), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I770 (.Y(N3208), .A0(N3714), .A1(N3808), .B0(N3625), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I771 (.Y(N3409), .A0(N3714), .A1(N4079), .B0(N3315), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I772 (.Y(N3621), .A(N3714), .B(N3522));
AOI22XL cynw_cm_float_rcp_I773 (.Y(N3292), .A0(N3714), .A1(N3489), .B0(N3724), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I774 (.Y(N3502), .A0(N3714), .A1(N4091), .B0(N3394), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I775 (.Y(N3706), .A0(N3714), .A1(a_man[16]), .B0(N3279), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I776 (.Y(N3908), .A0(N3714), .A1(N3488), .B0(N3419), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I777 (.Y(N4115), .A0(N3714), .A1(N3779), .B0(N4025), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I778 (.Y(N3381), .A0(N3714), .A1(N3811), .B0(N3506), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I779 (.Y(N3582), .A0(N3714), .A1(N4025), .B0(N3949), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I780 (.Y(N3788), .A0(N3714), .A1(N3693), .B0(N3913), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I781 (.Y(N3987), .A0(N3714), .A1(N3250), .B0(N3384), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I782 (.Y(N3955), .A0(N3714), .A1(N3825), .B0(N4102), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I783 (.Y(N3224), .A0(N3714), .A1(N3298), .B0(N3643), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I784 (.Y(N3428), .A0(N3714), .A1(N3590), .B0(N3779), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I785 (.Y(N3637), .A0(N3714), .A1(N3912), .B0(N3739), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I786 (.Y(N3839), .A0(N3714), .A1(N3761), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I787 (.Y(N4039), .A0(N3714), .A1(N3625), .B0(N4021), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I788 (.Y(N3313), .A0(N3714), .A1(N3586), .B0(N3795), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I789 (.Y(N3520), .A0(N3714), .A1(N3793), .B0(N3501), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I790 (.Y(N3721), .A0(N3714), .A1(N3990), .B0(N3910), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I791 (.Y(N3926), .A0(N3714), .A1(N3581), .B0(N3384), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I792 (.Y(N4129), .A0(N3714), .A1(N3269), .B0(N3581), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I793 (.Y(N3392), .A0(N3714), .A1(N3384), .B0(N3785), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I794 (.Y(N3599), .A0(N3714), .A1(N4078), .B0(N3985), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I795 (.Y(N3805), .A0(N3714), .A1(N3910), .B0(N3255), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I796 (.Y(N4002), .A0(N3714), .A1(N3550), .B0(N3260), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I797 (.Y(N3273), .A0(N3714), .A1(N4015), .B0(N3830), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I798 (.Y(N3480), .A0(N3714), .A1(N3958), .B0(N3399), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I799 (.Y(N3688), .A0(N3714), .A1(N4042), .B0(N3676), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I800 (.Y(N3887), .A0(N3714), .A1(N3431), .B0(N3399), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I801 (.Y(N4094), .A0(N3714), .A1(N3279), .B0(N4065), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I802 (.Y(N3363), .A0(N3714), .A1(N2381), .B0(N3452), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I803 (.Y(N3414), .A(N3752), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I804 (.Y(N3840), .A0(N3641), .A1(N3346), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I805 (.Y(N4026), .A0(N3641), .A1(N3465), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I806 (.Y(N4080), .A0(N3641), .A1(N3752), .B0(a_man[16]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I807 (.Y(N3551), .A(N3708));
AOI22XL cynw_cm_float_rcp_I808 (.Y(N3432), .A0(N3641), .A1(N4036), .B0(N3465), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I809 (.Y(N3974), .A0(N3641), .A1(a_man[16]), .B0(N3517), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I810 (.Y(N3660), .A0(N3641), .A1(N3344), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I811 (.Y(N3209), .A0(N3641), .A1(N3723), .B0(N3222), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I812 (.Y(N3295), .A(N3641), .B(N3869));
AOI22XL cynw_cm_float_rcp_I813 (.Y(N4117), .A0(N3641), .A1(N3517), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I814 (.Y(N3530), .A0(N3641), .A1(N3517), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I815 (.Y(N3317), .A0(N3641), .A1(N3465), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I816 (.Y(N3610), .A0(N3641), .A1(N3222), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I817 (.Y(N3248), .A0(N3641), .A1(N4036), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I818 (.Y(N3827), .A0(N3641), .A1(N3636), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I819 (.Y(N3299), .A0(N3641), .A1(N3482), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I820 (.Y(N3759), .A0(N3641), .A1(N3344), .B0(a_man[17]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I821 (.Y(N3960), .A(N3517));
NAND2XL cynw_cm_float_rcp_I822 (.Y(N3227), .A(N3344), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I823 (.Y(N4044), .A0(N3641), .A1(N4036), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I824 (.Y(N3319), .A0(N3641), .A1(N3636), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I825 (.Y(N3728), .A0(N3641), .A1(N3344), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I826 (.Y(N3931), .A0(N3641), .A1(N3752), .B0(N3482), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I827 (.Y(N3397), .A(a_man[18]), .B(N3346));
AOI22XL cynw_cm_float_rcp_I828 (.Y(N3726), .A0(N3641), .A1(N3222), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I829 (.Y(N3211), .A0(N3714), .A1(N3530), .B0(N3335), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I830 (.Y(N3412), .A0(N3714), .A1(N3384), .B0(N3414), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I831 (.Y(N3623), .A0(N3714), .A1(N3317), .B0(N3840), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I832 (.Y(N3824), .A0(N3714), .A1(N3570), .B0(N4026), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I833 (.Y(N4024), .A0(N3714), .A1(N3610), .B0(N3643), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I834 (.Y(N3297), .A0(N3714), .A1(N3390), .B0(N3643), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I835 (.Y(N3504), .A(N3643), .B(a_man[19]));
AOI22XL cynw_cm_float_rcp_I836 (.Y(N3259), .A0(N3714), .A1(N3808), .B0(N4080), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I837 (.Y(N3464), .A0(N3714), .A1(N3248), .B0(N3506), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I838 (.Y(N3675), .A0(N3714), .A1(N3739), .B0(N3551), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I839 (.Y(N3873), .A0(N3714), .A1(N3394), .B0(N3638), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I840 (.Y(N4077), .A0(N3714), .A1(N3739), .B0(N3860), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I841 (.Y(N3348), .A0(N3714), .A1(N3505), .B0(N3429), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I842 (.Y(N3549), .A0(N3714), .A1(N3548), .B0(N3432), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I843 (.Y(N3756), .A0(N3714), .A1(N3830), .B0(N3414), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I844 (.Y(N3956), .A(N3714), .B(N3827));
NOR2XL cynw_cm_float_rcp_I845 (.Y(N3430), .A(a_man[19]), .B(N3614));
AOI22XL cynw_cm_float_rcp_I846 (.Y(N4040), .A0(N3714), .A1(N3299), .B0(N3346), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I847 (.Y(N3316), .A0(N3714), .A1(N3570), .B0(N3395), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I848 (.Y(N3523), .A0(N3714), .A1(N4065), .B0(N3779), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I849 (.Y(N3725), .A0(N3714), .A1(N2381), .B0(N3666), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I850 (.Y(N3928), .A(a_man[19]), .B(N3384));
AOI22XL cynw_cm_float_rcp_I851 (.Y(N3483), .A0(N3714), .A1(N3335), .B0(N4073), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I852 (.Y(N3691), .A0(N3714), .A1(N3759), .B0(N3974), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I853 (.Y(N3888), .A0(N3714), .A1(N3960), .B0(N3641), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I854 (.Y(N4096), .A0(N3714), .A1(N3227), .B0(N3660), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I855 (.Y(N3366), .A0(N3714), .A1(N4003), .B0(N3976), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I856 (.Y(N3567), .A0(N3714), .A1(N3992), .B0(N3912), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I857 (.Y(N3772), .A0(N3714), .A1(N4044), .B0(N3785), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I858 (.Y(N3972), .A0(N3714), .A1(N3319), .B0(N3212), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I859 (.Y(N3241), .A0(N3714), .A1(N3958), .B0(N3949), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I860 (.Y(N3449), .A0(N3714), .A1(N3728), .B0(N3419), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I861 (.Y(N3656), .A0(N3714), .A1(N3931), .B0(N3209), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I862 (.Y(N3855), .A0(N3714), .A1(N3506), .B0(N3614), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I863 (.Y(N4057), .A0(N3714), .A1(N3397), .B0(N3672), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I864 (.Y(N3330), .A0(N3714), .A1(N3212), .B0(N3543), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I865 (.Y(N3537), .A0(N3714), .A1(N3298), .B0(N3761), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I866 (.Y(N3740), .A0(N3714), .A1(N3431), .B0(N3295), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I867 (.Y(N3939), .A0(N3714), .A1(N3676), .B0(N3469), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I868 (.Y(N3207), .A0(N3714), .A1(N3726), .B0(N4079), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I869 (.Y(N3408), .A0(N3714), .A1(N3958), .B0(N4117), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I870 (.Y(N3620), .A0(N3714), .A1(N4026), .B0(N3949), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I871 (.Y(N3822), .A0(N3714), .A1(N3643), .B0(N4137), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I872 (.Y(N4022), .A0(N3714), .A1(N3390), .B0(N4137), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I873 (.Y(N3786), .A0(N3411), .A1(N3211), .B0(N3889), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I874 (.Y(N3986), .A0(N3411), .A1(N3412), .B0(N4097), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I875 (.Y(N3256), .A0(N3411), .A1(N3623), .B0(N3367), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I876 (.Y(N3460), .A0(N3411), .A1(N3824), .B0(N3568), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I877 (.Y(N3670), .A0(N3411), .A1(N4024), .B0(N3854), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I878 (.Y(N3870), .A0(N3411), .A1(N3297), .B0(N3737), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I879 (.Y(N4071), .A(N3411), .B(N3504));
NOR2XL cynw_cm_float_rcp_I880 (.Y(N3798), .A(N3714), .B(N3390));
NOR2XL cynw_cm_float_rcp_I881 (.Y(N3954), .A(N3798), .B(a_man[20]));
AOI22XL cynw_cm_float_rcp_I882 (.Y(N4037), .A0(N3411), .A1(N3259), .B0(N3741), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I883 (.Y(N3311), .A0(N3411), .A1(N3464), .B0(N3942), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I884 (.Y(N3518), .A0(N3411), .A1(N3675), .B0(N3208), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I885 (.Y(N3719), .A0(N3411), .A1(N3873), .B0(N3409), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I886 (.Y(N3924), .A0(N3411), .A1(N4077), .B0(N3621), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I887 (.Y(N4127), .A0(N3411), .A1(N3348), .B0(N3292), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I888 (.Y(N3391), .A0(N3411), .A1(N3549), .B0(N3502), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I889 (.Y(N3597), .A0(N3411), .A1(N3756), .B0(N3706), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I890 (.Y(N3803), .A0(N3411), .A1(N3956), .B0(N3908), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I891 (.Y(N4000), .A0(N3411), .A1(N3430), .B0(N4115), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I892 (.Y(N3270), .A0(N3411), .A1(N4040), .B0(N3381), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I893 (.Y(N3478), .A0(N3411), .A1(N3316), .B0(N3582), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I894 (.Y(N3686), .A0(N3411), .A1(N3523), .B0(N3788), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I895 (.Y(N3885), .A0(N3411), .A1(N3725), .B0(N3987), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I896 (.Y(N4092), .A0(N3411), .A1(N3928), .B0(N3326), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I897 (.Y(N3651), .A0(N3411), .A1(N3483), .B0(N3955), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I898 (.Y(N3852), .A0(N3411), .A1(N3691), .B0(N3224), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I899 (.Y(N4052), .A0(N3411), .A1(N3888), .B0(N3428), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I900 (.Y(N3327), .A0(N3411), .A1(N4096), .B0(N3637), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I901 (.Y(N3533), .A0(N3411), .A1(N3366), .B0(N3839), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I902 (.Y(N3734), .A0(N3411), .A1(N3567), .B0(N4039), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I903 (.Y(N3937), .A0(N3411), .A1(N3772), .B0(N3313), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I904 (.Y(N3205), .A0(N3411), .A1(N3972), .B0(N3520), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I905 (.Y(N3405), .A0(N3411), .A1(N3241), .B0(N3721), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I906 (.Y(N3616), .A0(N3411), .A1(N3449), .B0(N3926), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I907 (.Y(N3818), .A0(N3411), .A1(N3656), .B0(N4129), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I908 (.Y(N4017), .A0(N3411), .A1(N3855), .B0(N3392), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I909 (.Y(N3287), .A0(N3411), .A1(N4057), .B0(N3599), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I910 (.Y(N3496), .A0(N3411), .A1(N3330), .B0(N3805), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I911 (.Y(N3699), .A0(N3411), .A1(N3537), .B0(N4002), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I912 (.Y(N3901), .A0(N3411), .A1(N3740), .B0(N3273), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I913 (.Y(N4109), .A0(N3411), .A1(N3939), .B0(N3480), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I914 (.Y(N3376), .A0(N3411), .A1(N3207), .B0(N3688), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I915 (.Y(N3576), .A0(N3411), .A1(N3408), .B0(N3887), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I916 (.Y(N3781), .A0(N3411), .A1(N3620), .B0(N4094), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I917 (.Y(N3981), .A0(N3411), .A1(N3822), .B0(N3363), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I918 (.Y(N3252), .A0(N3411), .A1(N4022), .B0(a_man[19]), .B1(a_man[20]));
OAI2BB1X1 cynw_cm_float_rcp_I919 (.Y(N3457), .A0N(N4137), .A1N(a_man[19]), .B0(N3411));
NOR2XL cynw_cm_float_rcp_I920 (.Y(N3358), .A(N3714), .B(N3452));
NOR2XL cynw_cm_float_rcp_I921 (.Y(N3866), .A(N3358), .B(a_man[20]));
INVX1 cynw_cm_float_rcp_I922 (.Y(N4114), .A(a_man[21]));
AOI22XL cynw_cm_float_rcp_I923 (.Y(N3218), .A0(N4114), .A1(N3786), .B0(N3820), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I924 (.Y(N3421), .A0(N4114), .A1(N3986), .B0(N4019), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I925 (.Y(N3631), .A0(N4114), .A1(N3256), .B0(N3290), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I926 (.Y(N3832), .A0(N4114), .A1(N3460), .B0(N3499), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I927 (.Y(N4029), .A0(N4114), .A1(N3670), .B0(N3702), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I928 (.Y(N3303), .A0(N4114), .A1(N3870), .B0(N3904), .B1(a_man[21]));
NAND2XL cynw_cm_float_rcp_I929 (.Y(N3510), .A(N4114), .B(N4071));
NOR2XL cynw_cm_float_rcp_I930 (.Y(N3917), .A(a_man[21]), .B(N4071));
NAND2XL cynw_cm_float_rcp_I931 (.Y(N3592), .A(N4114), .B(N3954));
AOI22XL cynw_cm_float_rcp_I932 (.Y(N3264), .A0(N4114), .A1(N4037), .B0(N4069), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I933 (.Y(N3471), .A0(N4114), .A1(N3311), .B0(N3341), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I934 (.Y(N3679), .A0(N4114), .A1(N3518), .B0(N3546), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I935 (.Y(N3878), .A0(N4114), .A1(N3719), .B0(N3749), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I936 (.Y(N4084), .A0(N4114), .A1(N3924), .B0(N3952), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I937 (.Y(N3354), .A0(N4114), .A1(N4127), .B0(N3220), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I938 (.Y(N3555), .A0(N4114), .A1(N3391), .B0(N3425), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I939 (.Y(N3763), .A0(N4114), .A1(N3597), .B0(N3634), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I940 (.Y(N3964), .A0(N4114), .A1(N3803), .B0(N3835), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I941 (.Y(N3231), .A0(N4114), .A1(N4000), .B0(N4033), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I942 (.Y(N3436), .A0(N4114), .A1(N3270), .B0(N3306), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I943 (.Y(N3645), .A0(N4114), .A1(N3478), .B0(N3513), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I944 (.Y(N3844), .A0(N4114), .A1(N3686), .B0(N3716), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I945 (.Y(N4048), .A0(N4114), .A1(N3885), .B0(N3920), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I946 (.Y(N3322), .A0(N4114), .A1(N4092), .B0(N4122), .B1(a_man[21]));
NOR2XL cynw_cm_float_rcp_I947 (.Y(N3848), .A(N3411), .B(N3711));
NOR2XL cynw_cm_float_rcp_I948 (.Y(N3528), .A(N3848), .B(a_man[21]));
AOI22XL cynw_cm_float_rcp_I949 (.Y(N3812), .A0(N4114), .A1(N3651), .B0(N3474), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I950 (.Y(N4009), .A0(N4114), .A1(N3852), .B0(N3682), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I951 (.Y(N3280), .A0(N4114), .A1(N4052), .B0(N3881), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I952 (.Y(N3490), .A0(N4114), .A1(N3327), .B0(N4087), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I953 (.Y(N3694), .A0(N4114), .A1(N3533), .B0(N3357), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I954 (.Y(N3894), .A0(N4114), .A1(N3734), .B0(N3558), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I955 (.Y(N4103), .A0(N4114), .A1(N3937), .B0(N3766), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I956 (.Y(N3371), .A0(N4114), .A1(N3205), .B0(N3967), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I957 (.Y(N3571), .A0(N4114), .A1(N3405), .B0(N3234), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I958 (.Y(N3776), .A0(N4114), .A1(N3616), .B0(N3439), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I959 (.Y(N3977), .A0(N4114), .A1(N3818), .B0(N3648), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I960 (.Y(N3246), .A0(N4114), .A1(N4017), .B0(N3847), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I961 (.Y(N3453), .A0(N4114), .A1(N3287), .B0(N4051), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I962 (.Y(N3662), .A0(N4114), .A1(N3496), .B0(N3325), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I963 (.Y(N3861), .A0(N4114), .A1(N3699), .B0(N3532), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I964 (.Y(N4062), .A0(N4114), .A1(N3901), .B0(N3732), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I965 (.Y(N3336), .A0(N4114), .A1(N4109), .B0(N3936), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I966 (.Y(N3540), .A0(N4114), .A1(N3376), .B0(N4136), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I967 (.Y(N3744), .A0(N4114), .A1(N3576), .B0(N3401), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I968 (.Y(N3945), .A0(N4114), .A1(N3781), .B0(N3612), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I969 (.Y(N3213), .A0(N4114), .A1(N3981), .B0(N3814), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I970 (.Y(N3415), .A0(N4114), .A1(N3252), .B0(N4012), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I971 (.Y(N3626), .A0(N4114), .A1(N3457), .B0(N3283), .B1(a_man[21]));
NAND2XL cynw_cm_float_rcp_I972 (.Y(N3826), .A(N4114), .B(N3866));
AOI22XL cynw_cm_float_rcp_I973 (.Y(N3618), .A0(N3641), .A1(N3346), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I974 (.Y(N3424), .A0(N3641), .A1(N3465), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I975 (.Y(N4032), .A0(N3641), .A1(N3636), .B0(N3723), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I976 (.Y(N3995), .A0(N3641), .A1(N3869), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I977 (.Y(N3943), .A0(N3641), .A1(N3708), .B0(N3465), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I978 (.Y(N3674), .A(N3723), .B(a_man[18]));
NOR2XL cynw_cm_float_rcp_I979 (.Y(N4076), .A(N3641), .B(N3346));
NAND2XL cynw_cm_float_rcp_I980 (.Y(N3755), .A(N3465), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I981 (.Y(N3771), .A0(N3641), .A1(N3869), .B0(N3222), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I982 (.Y(N3448), .A0(N3641), .A1(N3222), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I983 (.Y(N4056), .A0(N3641), .A1(a_man[17]), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I984 (.Y(N3751), .A0(N3714), .A1(N3384), .B0(N4117), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I985 (.Y(N3953), .A0(N3714), .A1(N3317), .B0(N3940), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I986 (.Y(N3221), .A0(N3714), .A1(N3923), .B0(N3494), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I987 (.Y(N3426), .A0(N3714), .A1(N3943), .B0(N3792), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I988 (.Y(N3635), .A0(N3714), .A1(N3209), .B0(N4065), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I989 (.Y(N3837), .A0(N3714), .A1(N4091), .B0(N4137), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I990 (.Y(N4035), .A0(N3714), .A1(N3384), .B0(N3452), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I991 (.Y(N3310), .A(N3714), .B(N2381));
AOI22XL cynw_cm_float_rcp_I992 (.Y(N3389), .A0(N3714), .A1(N3600), .B0(N3795), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I993 (.Y(N3595), .A0(N3714), .A1(N3586), .B0(N4134), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I994 (.Y(N3801), .A0(N3714), .A1(N3802), .B0(N3761), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I995 (.Y(N3998), .A0(N3714), .A1(N3394), .B0(N3840), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I996 (.Y(N3268), .A0(N3714), .A1(N3794), .B0(N3624), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I997 (.Y(N3477), .A0(N3714), .A1(N3794), .B0(N3522), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I998 (.Y(N3685), .A0(N3714), .A1(N3674), .B0(N3618), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I999 (.Y(N3884), .A0(N3714), .A1(N4076), .B0(N3384), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1000 (.Y(N4090), .A0(N3714), .A1(N3755), .B0(N3346), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1001 (.Y(N3360), .A0(N3714), .A1(N3840), .B0(N3395), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1002 (.Y(N3561), .A0(N3714), .A1(N3395), .B0(N3860), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1003 (.Y(N3768), .A0(N3714), .A1(N3976), .B0(N3830), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1004 (.Y(N3403), .A0(N3714), .A1(N3759), .B0(N3913), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1005 (.Y(N3613), .A0(N3714), .A1(N3940), .B0(N3469), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1006 (.Y(N3816), .A0(N3714), .A1(N3958), .B0(N3933), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1007 (.Y(N4014), .A0(N3714), .A1(N2381), .B0(N3618), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1008 (.Y(N3285), .A0(N3714), .A1(N3771), .B0(N3424), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1009 (.Y(N3493), .A0(N3714), .A1(a_man[18]), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1010 (.Y(N3697), .A0(N3714), .A1(N3448), .B0(N4032), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1011 (.Y(N3898), .A0(N3714), .A1(N3448), .B0(N3960), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1012 (.Y(N4106), .A0(N3714), .A1(N3976), .B0(N3242), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1013 (.Y(N3374), .A0(N3714), .A1(N4056), .B0(N3543), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1014 (.Y(N3574), .A0(N3714), .A1(N3641), .B0(N3969), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1015 (.Y(N3778), .A0(N3714), .A1(N3639), .B0(N3399), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1016 (.Y(N3979), .A0(N3714), .A1(N3494), .B0(N3526), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1017 (.Y(N3249), .A0(N3714), .A1(N3315), .B0(N3995), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1018 (.Y(N3455), .A0(N3714), .A1(N3891), .B0(N3260), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1019 (.Y(N3665), .A0(N3714), .A1(N3250), .B0(N3830), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1020 (.Y(N3864), .A(N3726), .B(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1021 (.Y(N3948), .A0(N3714), .A1(N3346), .B0(N3260), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1022 (.Y(N3216), .A0(N3714), .A1(a_man[17]), .B0(N3209), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1023 (.Y(N3418), .A0(N3714), .A1(N3535), .B0(N4091), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1024 (.Y(N3629), .A0(N3714), .A1(N2381), .B0(N3384), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I1025 (.Y(N3829), .A(N3714), .B(N2381));
NAND2XL cynw_cm_float_rcp_I1026 (.Y(N3332), .A(a_man[16]), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1027 (.Y(N3941), .A0(N3641), .A1(N3517), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1028 (.Y(N3907), .A0(N3641), .A1(N3723), .B0(N3344), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1029 (.Y(N3223), .A(N3641), .B(N3344));
AOI22XL cynw_cm_float_rcp_I1030 (.Y(N3838), .A0(N3641), .A1(N3222), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1031 (.Y(N3272), .A0(N3641), .A1(N3344), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1032 (.Y(N3362), .A0(N3641), .A1(N3344), .B0(N3222), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1033 (.Y(N3564), .A(N3641), .B(N3636));
AOI22XL cynw_cm_float_rcp_I1034 (.Y(N3237), .A0(N3641), .A1(N3869), .B0(N3482), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I1035 (.Y(N3444), .A(N3636), .B(a_man[18]));
NAND2XL cynw_cm_float_rcp_I1036 (.Y(N3605), .A(N3641), .B(N3636));
AOI22XL cynw_cm_float_rcp_I1037 (.Y(N4006), .A0(N3641), .A1(a_man[16]), .B0(N3723), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1038 (.Y(N3277), .A0(N3641), .A1(N3517), .B0(N3708), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1039 (.Y(N3485), .A(N3641), .B(N3482));
AOI22XL cynw_cm_float_rcp_I1040 (.Y(N4098), .A0(N3641), .A1(N3869), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1041 (.Y(N3791), .A0(N3641), .A1(N3723), .B0(N3517), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1042 (.Y(N4075), .A0(N3641), .A1(N3636), .B0(N3222), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1043 (.Y(N3225), .A0(N3641), .A1(N3344), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1044 (.Y(N3603), .A0(N3641), .A1(N3482), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1045 (.Y(N3275), .A0(N3641), .A1(N3869), .B0(N3752), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1046 (.Y(N3239), .A0(N3714), .A1(N3857), .B0(N3893), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1047 (.Y(N3446), .A0(N3714), .A1(N4026), .B0(N3550), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1048 (.Y(N3654), .A0(N3714), .A1(N3390), .B0(N4120), .B1(a_man[19]));
INVXL cynw_cm_float_rcp_I1049 (.Y(N3329), .A(N3488));
INVXL cynw_cm_float_rcp_I1050 (.Y(N3536), .A(N3301));
AOI22XL cynw_cm_float_rcp_I1051 (.Y(N3738), .A0(N3714), .A1(N3666), .B0(N3250), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1052 (.Y(N3703), .A0(N3714), .A1(N3605), .B0(N3332), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1053 (.Y(N3905), .A0(N3714), .A1(N4006), .B0(N3229), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1054 (.Y(N4112), .A0(N3714), .A1(N3277), .B0(N3941), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1055 (.Y(N3379), .A0(N3714), .A1(N3485), .B0(N3676), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1056 (.Y(N3578), .A0(N3714), .A1(N4098), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1057 (.Y(N3782), .A0(N3714), .A1(N3212), .B0(N3550), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1058 (.Y(N3983), .A0(N3714), .A1(N3958), .B0(N3466), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1059 (.Y(N3254), .A0(N3714), .A1(N3522), .B0(N3907), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1060 (.Y(N3459), .A0(N3714), .A1(N3223), .B0(N3876), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1061 (.Y(N3669), .A0(N3714), .A1(N4137), .B0(N3352), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1062 (.Y(N3868), .A0(N3714), .A1(N3452), .B0(N4101), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1063 (.Y(N4070), .A0(N3714), .A1(a_man[16]), .B0(N3808), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1064 (.Y(N3342), .A0(N3714), .A1(N3723), .B0(N3638), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1065 (.Y(N3750), .A0(N3714), .A1(N2381), .B0(N3643), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1066 (.Y(N3307), .A0(N3714), .A1(N3369), .B0(N3223), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1067 (.Y(N3514), .A0(N3714), .A1(N3791), .B0(N3838), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1068 (.Y(N3717), .A0(N3714), .A1(N3450), .B0(N3223), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1069 (.Y(N3921), .A0(N3714), .A1(N3625), .B0(N3317), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1070 (.Y(N4123), .A0(N3714), .A1(N4137), .B0(N3260), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1071 (.Y(N3387), .A0(N3714), .A1(N4075), .B0(N3279), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1072 (.Y(N3593), .A0(N3714), .A1(N3444), .B0(N3660), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1073 (.Y(N3799), .A0(N3714), .A1(N4117), .B0(N3856), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1074 (.Y(N3996), .A0(N3714), .A1(N3600), .B0(N3272), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1075 (.Y(N3266), .A0(N3714), .A1(N3225), .B0(N3242), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1076 (.Y(N3475), .A0(N3714), .A1(N3913), .B0(N3726), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1077 (.Y(N3683), .A0(N3714), .A1(N4091), .B0(N3362), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1078 (.Y(N3882), .A0(N3714), .A1(N3488), .B0(N3564), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1079 (.Y(N4088), .A0(N3714), .A1(N3793), .B0(N3237), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1080 (.Y(N3359), .A0(N3714), .A1(N3550), .B0(N3444), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1081 (.Y(N3559), .A0(N3714), .A1(N3444), .B0(N3260), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1082 (.Y(N3767), .A0(N3714), .A1(N3958), .B0(N3795), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1083 (.Y(N3968), .A0(N3714), .A1(N3603), .B0(a_man[18]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1084 (.Y(N3235), .A0(N3714), .A1(N3860), .B0(N3351), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1085 (.Y(N3440), .A0(N3714), .A1(N3526), .B0(N3876), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1086 (.Y(N3649), .A0(N3714), .A1(N3275), .B0(N3726), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1087 (.Y(N3849), .A0(N3714), .A1(N3641), .B0(N3643), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1088 (.Y(N3815), .A0(N3411), .A1(N3239), .B0(N3751), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1089 (.Y(N4013), .A0(N3411), .A1(N3446), .B0(N3953), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1090 (.Y(N3284), .A0(N3411), .A1(N3654), .B0(N3221), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1091 (.Y(N3492), .A0(N3411), .A1(N3346), .B0(N3426), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1092 (.Y(N3696), .A0(N3411), .A1(N3329), .B0(N3635), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1093 (.Y(N3897), .A0(N3411), .A1(N3536), .B0(N3837), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1094 (.Y(N4105), .A0(N3411), .A1(N3738), .B0(N4035), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1095 (.Y(N3373), .A0(N3411), .A1(N3711), .B0(N3310), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I1096 (.Y(N3573), .A(N3411), .B(N3711));
AOI22XL cynw_cm_float_rcp_I1097 (.Y(N3664), .A0(N3411), .A1(N3703), .B0(N3389), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1098 (.Y(N3863), .A0(N3411), .A1(N3905), .B0(N3595), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1099 (.Y(N4064), .A0(N3411), .A1(N4112), .B0(N3801), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1100 (.Y(N3338), .A0(N3411), .A1(N3379), .B0(N3998), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1101 (.Y(N3542), .A0(N3411), .A1(N3578), .B0(N3268), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1102 (.Y(N3746), .A0(N3411), .A1(N3782), .B0(N3477), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1103 (.Y(N3947), .A0(N3411), .A1(N3983), .B0(N3685), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1104 (.Y(N3215), .A0(N3411), .A1(N3254), .B0(N3884), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1105 (.Y(N3417), .A0(N3411), .A1(N3459), .B0(N4090), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1106 (.Y(N3628), .A0(N3411), .A1(N3669), .B0(N3360), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1107 (.Y(N3828), .A0(N3411), .A1(N3868), .B0(N3561), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1108 (.Y(N4027), .A0(N3411), .A1(N4070), .B0(N3768), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1109 (.Y(N3300), .A0(N3411), .A1(N3342), .B0(N3673), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1110 (.Y(N3508), .A0(N3411), .A1(N3447), .B0(N3872), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1111 (.Y(N3710), .A0(N3411), .A1(N3750), .B0(N3743), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1112 (.Y(N3915), .A0(N3411), .A1(N3928), .B0(N3743), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I1113 (.Y(N4119), .A(N3743), .B(a_man[20]));
NOR2XL cynw_cm_float_rcp_I1114 (.Y(N3589), .A(N3411), .B(N3560));
AOI22XL cynw_cm_float_rcp_I1115 (.Y(N3262), .A0(N3411), .A1(N3307), .B0(N3403), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1116 (.Y(N3468), .A0(N3411), .A1(N3514), .B0(N3613), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1117 (.Y(N3677), .A0(N3411), .A1(N3717), .B0(N3816), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1118 (.Y(N3875), .A0(N3411), .A1(N3921), .B0(N4014), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1119 (.Y(N4082), .A0(N3411), .A1(N4123), .B0(N3285), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1120 (.Y(N3350), .A0(N3411), .A1(N3387), .B0(N3493), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1121 (.Y(N3553), .A0(N3411), .A1(N3593), .B0(N3697), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1122 (.Y(N3760), .A0(N3411), .A1(N3799), .B0(N3898), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1123 (.Y(N3961), .A0(N3411), .A1(N3996), .B0(N4106), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1124 (.Y(N3228), .A0(N3411), .A1(N3266), .B0(N3374), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1125 (.Y(N3434), .A0(N3411), .A1(N3475), .B0(N3574), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1126 (.Y(N3642), .A0(N3411), .A1(N3683), .B0(N3778), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1127 (.Y(N3842), .A0(N3411), .A1(N3882), .B0(N3979), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1128 (.Y(N4045), .A0(N3411), .A1(N4088), .B0(N3249), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1129 (.Y(N3320), .A0(N3411), .A1(N3359), .B0(N3455), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1130 (.Y(N3525), .A0(N3411), .A1(N3559), .B0(N3665), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1131 (.Y(N3729), .A0(N3411), .A1(N3767), .B0(N3864), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1132 (.Y(N3932), .A0(N3411), .A1(N3968), .B0(N3538), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1133 (.Y(N4133), .A0(N3411), .A1(N3235), .B0(N3948), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1134 (.Y(N3398), .A0(N3411), .A1(N3440), .B0(N3216), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1135 (.Y(N3607), .A0(N3411), .A1(N3649), .B0(N3418), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1136 (.Y(N3809), .A0(N3411), .A1(N3849), .B0(N3629), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1137 (.Y(N4007), .A0(N3411), .A1(N3504), .B0(N3829), .B1(a_man[20]));
INVXL cynw_cm_float_rcp_I1138 (.Y(N4126), .A(N3752));
AOI22XL cynw_cm_float_rcp_I1139 (.Y(N3596), .A0(N3641), .A1(N3752), .B0(N3517), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1140 (.Y(N3999), .A0(N3641), .A1(a_man[17]), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1141 (.Y(N3733), .A0(N3641), .A1(a_man[17]), .B0(N3346), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1142 (.Y(N3404), .A0(N3641), .A1(a_man[16]), .B0(N3222), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1143 (.Y(N4108), .A0(N3641), .A1(N3344), .B0(N3708), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1144 (.Y(N4067), .A0(N3641), .A1(N3346), .B0(N3517), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1145 (.Y(N3293), .A0(N3641), .A1(N3517), .B0(N4036), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1146 (.Y(N4074), .A0(N3641), .A1(N4036), .B0(N3222), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1147 (.Y(N3601), .A0(N3641), .A1(N3636), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1148 (.Y(N3806), .A0(N3641), .A1(N3222), .B0(N3517), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1149 (.Y(N3289), .A0(N3714), .A1(N3992), .B0(N3319), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1150 (.Y(N3498), .A0(N3714), .A1(N3785), .B0(N4042), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1151 (.Y(N3701), .A0(N3714), .A1(N4046), .B0(N3431), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1152 (.Y(N3903), .A0(N3714), .A1(N3432), .B0(N3494), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1153 (.Y(N4111), .A0(N3714), .A1(N3419), .B0(N3992), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1154 (.Y(N3378), .A0(N3714), .A1(N4079), .B0(N3726), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1155 (.Y(N3577), .A0(N3714), .A1(N3693), .B0(N3390), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1156 (.Y(N3867), .A0(N3714), .A1(N4134), .B0(N4126), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1157 (.Y(N4068), .A0(N3714), .A1(N3494), .B0(N3590), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1158 (.Y(N3340), .A0(N3714), .A1(N3608), .B0(N3596), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1159 (.Y(N3545), .A0(N3714), .A1(N3293), .B0(N3610), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1160 (.Y(N3748), .A0(N3714), .A1(N4025), .B0(N3999), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1161 (.Y(N3951), .A0(N3714), .A1(N3608), .B0(N4044), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1162 (.Y(N3219), .A0(N3714), .A1(N3399), .B0(N3225), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1163 (.Y(N3423), .A0(N3714), .A1(N3397), .B0(N3548), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1164 (.Y(N3633), .A0(N3714), .A1(N3505), .B0(N3830), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1165 (.Y(N3834), .A0(N3714), .A1(N3299), .B0(N3827), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1166 (.Y(N4031), .A0(N3714), .A1(N3570), .B0(N3614), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1167 (.Y(N3305), .A0(N3714), .A1(N3494), .B0(N3317), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1168 (.Y(N3512), .A0(N3714), .A1(N3399), .B0(N3759), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1169 (.Y(N3715), .A0(N3714), .A1(N4074), .B0(N3614), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1170 (.Y(N3919), .A0(N3714), .A1(N3641), .B0(N3384), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1171 (.Y(N3473), .A0(N3714), .A1(N3299), .B0(N3733), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1172 (.Y(N3681), .A0(N3714), .A1(N3913), .B0(N3899), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1173 (.Y(N3880), .A0(N3714), .A1(N3248), .B0(N3913), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1174 (.Y(N4086), .A0(N3714), .A1(N3399), .B0(N3404), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1175 (.Y(N3356), .A0(N3714), .A1(N3431), .B0(N3724), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1176 (.Y(N3557), .A0(N3714), .A1(N4074), .B0(N3419), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1177 (.Y(N3765), .A0(N3714), .A1(N3860), .B0(N3625), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1178 (.Y(N3966), .A0(N3714), .A1(N3601), .B0(N4079), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1179 (.Y(N3233), .A0(N3714), .A1(N3806), .B0(N3269), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1180 (.Y(N3438), .A0(N3714), .A1(N3601), .B0(N4108), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1181 (.Y(N3647), .A0(N3714), .A1(N3840), .B0(N3811), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1182 (.Y(N3846), .A0(N3714), .A1(N3448), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1183 (.Y(N4050), .A0(N3714), .A1(N3227), .B0(N3899), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1184 (.Y(N3324), .A0(N3714), .A1(N4102), .B0(N3857), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1185 (.Y(N3531), .A0(N3714), .A1(N4108), .B0(N3674), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1186 (.Y(N3731), .A0(N3714), .A1(N4044), .B0(N4067), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1187 (.Y(N3935), .A0(N3714), .A1(N3771), .B0(N3929), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1188 (.Y(N4135), .A0(N3714), .A1(N3346), .B0(N3494), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1189 (.Y(N3400), .A0(N3714), .A1(N3488), .B0(N3526), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1190 (.Y(N3611), .A0(N3714), .A1(N3212), .B0(N3494), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1191 (.Y(N4011), .A0(N3714), .A1(N3384), .B0(N4120), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1192 (.Y(N3282), .A0(N3714), .A1(N3384), .B0(N4015), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1193 (.Y(N3276), .A(N3222), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1194 (.Y(N4055), .A0(N3641), .A1(N3517), .B0(N3723), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1195 (.Y(N3580), .A0(N3641), .A1(N3708), .B0(N3869), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1196 (.Y(N3784), .A0(N3641), .A1(N3344), .B0(N3346), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1197 (.Y(N3343), .A(a_man[18]), .B(N3708));
AOI22XL cynw_cm_float_rcp_I1198 (.Y(N3309), .A0(N3641), .A1(N3869), .B0(N3465), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I1199 (.Y(N3516), .A(N3641), .B(N3482));
AOI22XL cynw_cm_float_rcp_I1200 (.Y(N4125), .A0(N3641), .A1(N3346), .B0(N3723), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I1201 (.Y(N3413), .A(N4036));
NAND2XL cynw_cm_float_rcp_I1202 (.Y(N3911), .A(N3482), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1203 (.Y(N3657), .A0(N3641), .A1(N3222), .B0(N3636), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1204 (.Y(N3331), .A0(N3641), .A1(N3222), .B0(N3482), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1205 (.Y(N3257), .A0(N3714), .A1(N3724), .B0(N3562), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1206 (.Y(N3461), .A0(N3714), .A1(N4102), .B0(N4067), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1207 (.Y(N3671), .A0(N3714), .A1(N3933), .B0(N3825), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1208 (.Y(N3871), .A0(N3714), .A1(N3526), .B0(N3390), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1209 (.Y(N4072), .A0(N3714), .A1(N3992), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1210 (.Y(N3345), .A0(N3714), .A1(N3494), .B0(N3488), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1211 (.Y(N3547), .A0(N3714), .A1(N3229), .B0(N3779), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1212 (.Y(N3753), .A0(N3714), .A1(N4015), .B0(N4137), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1213 (.Y(N4038), .A0(N3714), .A1(N3413), .B0(N3985), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1214 (.Y(N3312), .A0(N3714), .A1(N3992), .B0(N3276), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1215 (.Y(N3519), .A0(N3714), .A1(N4099), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1216 (.Y(N3720), .A0(N3714), .A1(N3580), .B0(N3332), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1217 (.Y(N3925), .A0(N3714), .A1(N3596), .B0(N3969), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1218 (.Y(N4128), .A(N3714), .B(N3995));
AOI22XL cynw_cm_float_rcp_I1219 (.Y(N3598), .A0(N3714), .A1(N3530), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1220 (.Y(N3804), .A0(N3714), .A1(N3911), .B0(N3754), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1221 (.Y(N4001), .A0(N3714), .A1(N3689), .B0(N4055), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1222 (.Y(N3271), .A0(N3714), .A1(N3933), .B0(N3923), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1223 (.Y(N3479), .A0(N3714), .A1(N3755), .B0(N3625), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1224 (.Y(N3687), .A0(N3714), .A1(N4073), .B0(N3723), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1225 (.Y(N3886), .A0(N3714), .A1(N3840), .B0(N3469), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1226 (.Y(N4093), .A0(N3714), .A1(a_man[17]), .B0(N4025), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1227 (.Y(N3361), .A0(N3714), .A1(a_man[18]), .B0(N3693), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1228 (.Y(N3563), .A(N3666), .B(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1229 (.Y(N3443), .A0(N3714), .A1(N3676), .B0(N3733), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1230 (.Y(N3652), .A0(N3714), .A1(N3564), .B0(N4065), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1231 (.Y(N3853), .A0(N3714), .A1(N3565), .B0(N3580), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1232 (.Y(N4053), .A0(N3714), .A1(N3424), .B0(N3784), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1233 (.Y(N3328), .A0(N3714), .A1(N4080), .B0(N3351), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1234 (.Y(N3534), .A0(N3714), .A1(N3309), .B0(N4108), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1235 (.Y(N3735), .A0(N3714), .A1(N4046), .B0(N3352), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1236 (.Y(N3938), .A0(N3714), .A1(N3601), .B0(N3643), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1237 (.Y(N3206), .A0(N3714), .A1(N4056), .B0(N3610), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1238 (.Y(N3406), .A0(N3714), .A1(N3674), .B0(N3343), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1239 (.Y(N3617), .A0(N3714), .A1(N3856), .B0(N3874), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1240 (.Y(N3819), .A0(N3714), .A1(N4058), .B0(N3899), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1241 (.Y(N4018), .A0(N3714), .A1(N3657), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1242 (.Y(N3288), .A0(N3714), .A1(N3301), .B0(N3309), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1243 (.Y(N3497), .A0(N3714), .A1(N3352), .B0(N3516), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1244 (.Y(N3700), .A0(N3714), .A1(N3331), .B0(N3838), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1245 (.Y(N3902), .A0(N3714), .A1(N3564), .B0(N4125), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1246 (.Y(N4110), .A0(N3714), .A1(N4120), .B0(N3787), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I1247 (.Y(N3377), .A(N3714), .B(N3335));
AOI22XL cynw_cm_float_rcp_I1248 (.Y(N3982), .A0(N3714), .A1(N3346), .B0(N3840), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1249 (.Y(N3253), .A0(N3714), .A1(N3723), .B0(N3603), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1250 (.Y(N3458), .A0(N3714), .A1(N3641), .B0(N3301), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I1251 (.Y(N3668), .A(N3714), .B(N3250));
AOI22XL cynw_cm_float_rcp_I1252 (.Y(N3422), .A0(N3411), .A1(N3257), .B0(N3289), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1253 (.Y(N3632), .A0(N3411), .A1(N3461), .B0(N3498), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1254 (.Y(N3833), .A0(N3411), .A1(N3671), .B0(N3701), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1255 (.Y(N4030), .A0(N3411), .A1(N3871), .B0(N3903), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1256 (.Y(N3304), .A0(N3411), .A1(N4072), .B0(N4111), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1257 (.Y(N3511), .A0(N3411), .A1(N3345), .B0(N3378), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1258 (.Y(N3713), .A0(N3411), .A1(N3547), .B0(N3577), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1259 (.Y(N3918), .A0(N3411), .A1(N3753), .B0(N3655), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1260 (.Y(N3994), .A0(N3411), .A1(N4038), .B0(N3867), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1261 (.Y(N3265), .A0(N3411), .A1(N3312), .B0(N4068), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1262 (.Y(N3472), .A0(N3411), .A1(N3519), .B0(N3340), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1263 (.Y(N3680), .A0(N3411), .A1(N3720), .B0(N3545), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1264 (.Y(N3879), .A0(N3411), .A1(N3925), .B0(N3748), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1265 (.Y(N4085), .A0(N3411), .A1(N4128), .B0(N3951), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1266 (.Y(N3355), .A0(N3411), .A1(N3598), .B0(N3219), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1267 (.Y(N3556), .A0(N3411), .A1(N3804), .B0(N3423), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1268 (.Y(N3764), .A0(N3411), .A1(N4001), .B0(N3633), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1269 (.Y(N3965), .A0(N3411), .A1(N3271), .B0(N3834), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1270 (.Y(N3232), .A0(N3411), .A1(N3479), .B0(N4031), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1271 (.Y(N3437), .A0(N3411), .A1(N3687), .B0(N3305), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1272 (.Y(N3646), .A0(N3411), .A1(N3886), .B0(N3512), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1273 (.Y(N3845), .A0(N3411), .A1(N4093), .B0(N3715), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1274 (.Y(N4049), .A0(N3411), .A1(N3361), .B0(N3919), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1275 (.Y(N3323), .A0(N3411), .A1(N3563), .B0(N3737), .B1(a_man[20]));
NOR2XL cynw_cm_float_rcp_I1276 (.Y(N3529), .A(N3411), .B(N4054));
AOI22XL cynw_cm_float_rcp_I1277 (.Y(N3609), .A0(N3411), .A1(N3443), .B0(N3473), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1278 (.Y(N3813), .A0(N3411), .A1(N3652), .B0(N3681), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1279 (.Y(N4010), .A0(N3411), .A1(N3853), .B0(N3880), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1280 (.Y(N3281), .A0(N3411), .A1(N4053), .B0(N4086), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1281 (.Y(N3491), .A0(N3411), .A1(N3328), .B0(N3356), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1282 (.Y(N3695), .A0(N3411), .A1(N3534), .B0(N3557), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1283 (.Y(N3895), .A0(N3411), .A1(N3735), .B0(N3765), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1284 (.Y(N4104), .A0(N3411), .A1(N3938), .B0(N3966), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1285 (.Y(N3372), .A0(N3411), .A1(N3206), .B0(N3233), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1286 (.Y(N3572), .A0(N3411), .A1(N3406), .B0(N3438), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1287 (.Y(N3777), .A0(N3411), .A1(N3617), .B0(N3647), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1288 (.Y(N3978), .A0(N3411), .A1(N3819), .B0(N3846), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1289 (.Y(N3247), .A0(N3411), .A1(N4018), .B0(N4050), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1290 (.Y(N3454), .A0(N3411), .A1(N3288), .B0(N3324), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1291 (.Y(N3663), .A0(N3411), .A1(N3497), .B0(N3531), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1292 (.Y(N3862), .A0(N3411), .A1(N3700), .B0(N3731), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1293 (.Y(N4063), .A0(N3411), .A1(N3902), .B0(N3935), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1294 (.Y(N3337), .A0(N3411), .A1(N4110), .B0(N4135), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1295 (.Y(N3541), .A0(N3411), .A1(N3377), .B0(N3400), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1296 (.Y(N3745), .A0(N3411), .A1(N3982), .B0(N3611), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1297 (.Y(N3946), .A0(N3411), .A1(N3253), .B0(N3673), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1298 (.Y(N3214), .A0(N3411), .A1(N3458), .B0(N4011), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1299 (.Y(N3416), .A0(N3411), .A1(N3668), .B0(N3282), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I1300 (.Y(N3627), .A(N3310), .B(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1301 (.Y(N3507), .A0(N4114), .A1(N3422), .B0(N3815), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1302 (.Y(N3709), .A0(N4114), .A1(N3632), .B0(N4013), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1303 (.Y(N3914), .A0(N4114), .A1(N3833), .B0(N3284), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1304 (.Y(N4118), .A0(N4114), .A1(N4030), .B0(N3492), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1305 (.Y(N3385), .A0(N4114), .A1(N3304), .B0(N3696), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1306 (.Y(N3588), .A0(N4114), .A1(N3511), .B0(N3897), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1307 (.Y(N3796), .A0(N4114), .A1(N3713), .B0(N4105), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1308 (.Y(N3991), .A0(N4114), .A1(N3918), .B0(N3373), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1309 (.Y(N3261), .A0(N4114), .A1(N3866), .B0(N3573), .B1(a_man[21]));
NOR2XL cynw_cm_float_rcp_I1310 (.Y(N3402), .A(a_man[20]), .B(N3326));
NOR2XL cynw_cm_float_rcp_I1311 (.Y(N3467), .A(N3402), .B(N4114));
AOI22XL cynw_cm_float_rcp_I1312 (.Y(N4081), .A0(N4114), .A1(N3994), .B0(N3664), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1313 (.Y(N3349), .A0(N4114), .A1(N3265), .B0(N3863), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1314 (.Y(N3552), .A0(N4114), .A1(N3472), .B0(N4064), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1315 (.Y(N3758), .A0(N4114), .A1(N3680), .B0(N3338), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1316 (.Y(N3959), .A0(N4114), .A1(N3879), .B0(N3542), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1317 (.Y(N3226), .A0(N4114), .A1(N4085), .B0(N3746), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1318 (.Y(N3433), .A0(N4114), .A1(N3355), .B0(N3947), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1319 (.Y(N3640), .A0(N4114), .A1(N3556), .B0(N3215), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1320 (.Y(N3841), .A0(N4114), .A1(N3764), .B0(N3417), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1321 (.Y(N4043), .A0(N4114), .A1(N3965), .B0(N3628), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1322 (.Y(N3318), .A0(N4114), .A1(N3232), .B0(N3828), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1323 (.Y(N3524), .A0(N4114), .A1(N3437), .B0(N4027), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1324 (.Y(N3727), .A0(N4114), .A1(N3646), .B0(N3300), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1325 (.Y(N3930), .A0(N4114), .A1(N3845), .B0(N3508), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1326 (.Y(N4132), .A0(N4114), .A1(N4049), .B0(N3710), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1327 (.Y(N3396), .A0(N4114), .A1(N3323), .B0(N3915), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1328 (.Y(N3606), .A0(N4114), .A1(N3529), .B0(N4119), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1329 (.Y(N3278), .A0(N4114), .A1(N3609), .B0(N3262), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1330 (.Y(N3487), .A0(N4114), .A1(N3813), .B0(N3468), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1331 (.Y(N3692), .A0(N4114), .A1(N4010), .B0(N3677), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1332 (.Y(N3892), .A0(N4114), .A1(N3281), .B0(N3875), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1333 (.Y(N4100), .A0(N4114), .A1(N3491), .B0(N4082), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1334 (.Y(N3370), .A0(N4114), .A1(N3695), .B0(N3350), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1335 (.Y(N3569), .A0(N4114), .A1(N3895), .B0(N3553), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1336 (.Y(N3775), .A0(N4114), .A1(N4104), .B0(N3760), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1337 (.Y(N3975), .A0(N4114), .A1(N3372), .B0(N3961), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1338 (.Y(N3245), .A0(N4114), .A1(N3572), .B0(N3228), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1339 (.Y(N3451), .A0(N4114), .A1(N3777), .B0(N3434), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1340 (.Y(N3661), .A0(N4114), .A1(N3978), .B0(N3642), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1341 (.Y(N3859), .A0(N4114), .A1(N3247), .B0(N3842), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1342 (.Y(N4061), .A0(N4114), .A1(N3454), .B0(N4045), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1343 (.Y(N3334), .A0(N4114), .A1(N3663), .B0(N3320), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1344 (.Y(N3539), .A0(N4114), .A1(N3862), .B0(N3525), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1345 (.Y(N3742), .A0(N4114), .A1(N4063), .B0(N3729), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1346 (.Y(N3944), .A0(N4114), .A1(N3337), .B0(N3932), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1347 (.Y(N3210), .A0(N4114), .A1(N3541), .B0(N4133), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1348 (.Y(N3410), .A0(N4114), .A1(N3745), .B0(N3398), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1349 (.Y(N3622), .A0(N4114), .A1(N3946), .B0(N3607), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1350 (.Y(N3823), .A0(N4114), .A1(N3214), .B0(N3809), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1351 (.Y(N4023), .A0(N4114), .A1(N3416), .B0(N4007), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1352 (.Y(N3296), .A0(N4114), .A1(N3627), .B0(N4071), .B1(a_man[21]));
INVX1 cynw_cm_float_rcp_I1353 (.Y(N3427), .A(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1354 (.Y(N449), .A0(N3427), .A1(N3507), .B0(N3218), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1355 (.Y(N450), .A0(N3427), .A1(N3709), .B0(N3421), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1356 (.Y(N451), .A0(N3427), .A1(N3914), .B0(N3631), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1357 (.Y(N452), .A0(N3427), .A1(N4118), .B0(N3832), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1358 (.Y(N453), .A0(N3427), .A1(N3385), .B0(N4029), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1359 (.Y(N454), .A0(N3427), .A1(N3588), .B0(N3303), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1360 (.Y(N455), .A0(N3427), .A1(N3796), .B0(N3510), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1361 (.Y(N456), .A0(N3427), .A1(N3991), .B0(N3917), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1362 (.Y(N457), .A0(N3427), .A1(N3261), .B0(N3592), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1364 (.Y(inst_cellmath__51[0]), .A0(N3427), .A1(N4081), .B0(N3264), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1365 (.Y(inst_cellmath__51[1]), .A0(N3427), .A1(N3349), .B0(N3471), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1366 (.Y(inst_cellmath__51[2]), .A0(N3427), .A1(N3552), .B0(N3679), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1367 (.Y(inst_cellmath__51[3]), .A0(N3427), .A1(N3758), .B0(N3878), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1368 (.Y(inst_cellmath__51[4]), .A0(N3427), .A1(N3959), .B0(N4084), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1369 (.Y(inst_cellmath__51[5]), .A0(N3427), .A1(N3226), .B0(N3354), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1370 (.Y(inst_cellmath__51[6]), .A0(N3427), .A1(N3433), .B0(N3555), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1371 (.Y(inst_cellmath__51[7]), .A0(N3427), .A1(N3640), .B0(N3763), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1372 (.Y(inst_cellmath__51[8]), .A0(N3427), .A1(N3841), .B0(N3964), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1373 (.Y(inst_cellmath__51[9]), .A0(N3427), .A1(N4043), .B0(N3231), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1374 (.Y(inst_cellmath__51[10]), .A0(N3427), .A1(N3318), .B0(N3436), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1375 (.Y(inst_cellmath__51[11]), .A0(N3427), .A1(N3524), .B0(N3645), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1376 (.Y(inst_cellmath__51[12]), .A0(N3427), .A1(N3727), .B0(N3844), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1377 (.Y(inst_cellmath__51[13]), .A0(N3427), .A1(N3930), .B0(N4048), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1378 (.Y(inst_cellmath__51[14]), .A0(N3427), .A1(N4132), .B0(N3322), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1379 (.Y(inst_cellmath__51[15]), .A0(N3427), .A1(N3396), .B0(N3528), .B1(a_man[22]));
NOR2XL cynw_cm_float_rcp_I1380 (.Y(inst_cellmath__51[16]), .A(a_man[22]), .B(N3606));
OAI2BB1X1 cynw_cm_float_rcp_I1381 (.Y(inst_cellmath__51[17]), .A0N(N3589), .A1N(a_man[21]), .B0(N3427));
AOI22XL cynw_cm_float_rcp_I1382 (.Y(N477), .A0(N3427), .A1(N3278), .B0(N3812), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1383 (.Y(N478), .A0(N3427), .A1(N3487), .B0(N4009), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1384 (.Y(N479), .A0(N3427), .A1(N3692), .B0(N3280), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1385 (.Y(N480), .A0(N3427), .A1(N3892), .B0(N3490), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1386 (.Y(N481), .A0(N3427), .A1(N4100), .B0(N3694), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1387 (.Y(N482), .A0(N3427), .A1(N3370), .B0(N3894), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1388 (.Y(N483), .A0(N3427), .A1(N3569), .B0(N4103), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1389 (.Y(N484), .A0(N3427), .A1(N3775), .B0(N3371), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1390 (.Y(N485), .A0(N3427), .A1(N3975), .B0(N3571), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1391 (.Y(N486), .A0(N3427), .A1(N3245), .B0(N3776), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1392 (.Y(N487), .A0(N3427), .A1(N3451), .B0(N3977), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1393 (.Y(N488), .A0(N3427), .A1(N3661), .B0(N3246), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1394 (.Y(N489), .A0(N3427), .A1(N3859), .B0(N3453), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1395 (.Y(N490), .A0(N3427), .A1(N4061), .B0(N3662), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1396 (.Y(N491), .A0(N3427), .A1(N3334), .B0(N3861), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1397 (.Y(N492), .A0(N3427), .A1(N3539), .B0(N4062), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1398 (.Y(N493), .A0(N3427), .A1(N3742), .B0(N3336), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1399 (.Y(N494), .A0(N3427), .A1(N3944), .B0(N3540), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1400 (.Y(N495), .A0(N3427), .A1(N3210), .B0(N3744), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1401 (.Y(N496), .A0(N3427), .A1(N3410), .B0(N3945), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1402 (.Y(N497), .A0(N3427), .A1(N3622), .B0(N3213), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1403 (.Y(N498), .A0(N3427), .A1(N3823), .B0(N3415), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1404 (.Y(N499), .A0(N3427), .A1(N4023), .B0(N3626), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1405 (.Y(N500), .A0(N3427), .A1(N3296), .B0(N3826), .B1(a_man[22]));
NOR2XL cynw_cm_float_rcp_I1406 (.Y(N3896), .A(N4114), .B(N3954));
XOR2XL inst_cellmath__62_0_I5051 (.Y(N5382), .A(N2871), .B(N2652));
XOR2XL inst_cellmath__62_0_I5052 (.Y(N5117), .A(N2749), .B(N2795));
XOR2XL inst_cellmath__62_0_I5053 (.Y(N5188), .A(N2766), .B(N2610));
XOR2XL inst_cellmath__62_0_I5054 (.Y(N5261), .A(N2603), .B(N2752));
XOR2XL inst_cellmath__62_0_I5055 (.Y(N5336), .A(N2580), .B(N2893));
XOR2XL inst_cellmath__62_0_I5056 (.Y(N5074), .A(N2690), .B(N2710));
XOR2XL inst_cellmath__62_0_I5057 (.Y(N5148), .A(N2627), .B(N2852));
XOR2XL inst_cellmath__62_0_I5058 (.Y(N5221), .A(N2703), .B(N2667));
INVX2 inst_cellmath__62_0_I1416 (.Y(N5294), .A(inst_cellmath__60[21]));
INVX2 inst_cellmath__62_0_I1417 (.Y(N5367), .A(inst_cellmath__60[22]));
BUFX3 inst_cellmath__62_0_I5061 (.Y(N11739), .A(inst_cellmath__60[23]));
INVX2 inst_cellmath__62_0_I1419 (.Y(N5176), .A(inst_cellmath__60[24]));
INVXL inst_cellmath__62_0_I1420 (.Y(N5248), .A(N449));
NOR2XL inst_cellmath__62_0_I1421 (.Y(inst_cellmath__62__W0[4]), .A(N5248), .B(N5382));
NOR2XL inst_cellmath__62_0_I1422 (.Y(inst_cellmath__62__W1[5]), .A(N5248), .B(N5117));
NOR2XL inst_cellmath__62_0_I1423 (.Y(N5158), .A(N5248), .B(N5188));
NOR2XL inst_cellmath__62_0_I1424 (.Y(N5302), .A(N5248), .B(N5261));
NOR2XL inst_cellmath__62_0_I1425 (.Y(N5112), .A(N5248), .B(N5336));
NOR2XL inst_cellmath__62_0_I1426 (.Y(N5258), .A(N5248), .B(N5074));
NOR2XL inst_cellmath__62_0_I1427 (.Y(N5069), .A(N5248), .B(N5148));
NOR2XL inst_cellmath__62_0_I1428 (.Y(N5216), .A(N5248), .B(N5221));
NOR2X2 inst_cellmath__62_0_I1429 (.Y(N5365), .A(N5248), .B(N5294));
NOR2X1 inst_cellmath__62_0_I1430 (.Y(N5174), .A(N5248), .B(N5367));
NOR2X2 inst_cellmath__62_0_I1431 (.Y(N5320), .A(N5248), .B(N11739));
NOR2XL inst_cellmath__62_0_I1432 (.Y(N5129), .A(N5248), .B(N5176));
INVXL inst_cellmath__62_0_I1433 (.Y(N5324), .A(N450));
NOR2XL inst_cellmath__62_0_I1434 (.Y(inst_cellmath__62__W0[5]), .A(N5324), .B(N5382));
NOR2XL inst_cellmath__62_0_I1435 (.Y(inst_cellmath__62__W0[6]), .A(N5324), .B(N5117));
NOR2XL inst_cellmath__62_0_I1436 (.Y(N5369), .A(N5324), .B(N5188));
NOR2XL inst_cellmath__62_0_I1437 (.Y(N5178), .A(N5324), .B(N5261));
NOR2XL inst_cellmath__62_0_I1438 (.Y(N5327), .A(N5324), .B(N5336));
NOR2XL inst_cellmath__62_0_I1439 (.Y(N5136), .A(N5324), .B(N5074));
NOR2XL inst_cellmath__62_0_I1440 (.Y(N5282), .A(N5324), .B(N5148));
NOR2XL inst_cellmath__62_0_I1441 (.Y(N5091), .A(N5324), .B(N5221));
NOR2XL inst_cellmath__62_0_I1442 (.Y(N5238), .A(N5324), .B(N5294));
NOR2XL inst_cellmath__62_0_I1443 (.Y(N5388), .A(N5324), .B(N5367));
NOR2XL inst_cellmath__62_0_I1444 (.Y(N5197), .A(N5324), .B(inst_cellmath__60[23]));
NOR2X1 inst_cellmath__62_0_I1445 (.Y(N5342), .A(N5324), .B(N5176));
INVXL inst_cellmath__62_0_I1446 (.Y(N5399), .A(N451));
NOR2XL inst_cellmath__62_0_I1447 (.Y(N5289), .A(N5399), .B(N5382));
NOR2XL inst_cellmath__62_0_I1448 (.Y(N5097), .A(N5399), .B(N5117));
NOR2XL inst_cellmath__62_0_I1449 (.Y(N5243), .A(N5399), .B(N5188));
NOR2XL inst_cellmath__62_0_I1450 (.Y(N5393), .A(N5399), .B(N5261));
NOR2XL inst_cellmath__62_0_I1451 (.Y(N5201), .A(N5399), .B(N5336));
NOR2XL inst_cellmath__62_0_I1452 (.Y(N5348), .A(N5399), .B(N5074));
NOR2XL inst_cellmath__62_0_I1453 (.Y(N5160), .A(N5399), .B(N5148));
NOR2XL inst_cellmath__62_0_I1454 (.Y(N5306), .A(N5399), .B(N5221));
NOR2XL inst_cellmath__62_0_I1455 (.Y(N5116), .A(N5399), .B(N5294));
NOR2XL inst_cellmath__62_0_I1456 (.Y(N5262), .A(N5399), .B(N5367));
NOR2XL inst_cellmath__62_0_I1457 (.Y(N5073), .A(N5399), .B(N11739));
NOR2X2 inst_cellmath__62_0_I1458 (.Y(N5220), .A(N5399), .B(N5176));
INVXL inst_cellmath__62_0_I1459 (.Y(N5134), .A(N452));
NOR2XL inst_cellmath__62_0_I1460 (.Y(N5165), .A(N5134), .B(N5382));
NOR2XL inst_cellmath__62_0_I1461 (.Y(N5311), .A(N5134), .B(N5117));
NOR2XL inst_cellmath__62_0_I1462 (.Y(N5122), .A(N5134), .B(N5188));
NOR2XL inst_cellmath__62_0_I1463 (.Y(N5267), .A(N5134), .B(N5261));
NOR2XL inst_cellmath__62_0_I1464 (.Y(N5078), .A(N5134), .B(N5336));
NOR2XL inst_cellmath__62_0_I1465 (.Y(N5226), .A(N5134), .B(N5074));
NOR2XL inst_cellmath__62_0_I1466 (.Y(N5374), .A(N5134), .B(N5148));
NOR2XL inst_cellmath__62_0_I1467 (.Y(N5181), .A(N5134), .B(N5221));
NOR2XL inst_cellmath__62_0_I1468 (.Y(N5330), .A(N5134), .B(N5294));
NOR2XL inst_cellmath__62_0_I1469 (.Y(N5141), .A(N5134), .B(N5367));
NOR2XL inst_cellmath__62_0_I1470 (.Y(N5286), .A(N5134), .B(N11739));
NOR2XL inst_cellmath__62_0_I1471 (.Y(N5094), .A(N5134), .B(N5176));
INVXL inst_cellmath__62_0_I1472 (.Y(N5207), .A(N453));
NOR2XL inst_cellmath__62_0_I1473 (.Y(N5381), .A(N5207), .B(N5382));
NOR2XL inst_cellmath__62_0_I1474 (.Y(N5187), .A(N5207), .B(N5117));
NOR2XL inst_cellmath__62_0_I1475 (.Y(N5335), .A(N5207), .B(N5188));
NOR2XL inst_cellmath__62_0_I1476 (.Y(N5147), .A(N5207), .B(N5261));
NOR2XL inst_cellmath__62_0_I1477 (.Y(N5293), .A(N5207), .B(N5336));
NOR2XL inst_cellmath__62_0_I1478 (.Y(N5101), .A(N5207), .B(N5074));
NOR2XL inst_cellmath__62_0_I1479 (.Y(N5247), .A(N5207), .B(N5148));
NOR2XL inst_cellmath__62_0_I1480 (.Y(N5398), .A(N5207), .B(N5221));
NOR2XL inst_cellmath__62_0_I1481 (.Y(N5206), .A(N5207), .B(N5294));
NOR2XL inst_cellmath__62_0_I1482 (.Y(N5355), .A(N5207), .B(N5367));
NOR2XL inst_cellmath__62_0_I1483 (.Y(N5164), .A(N5207), .B(N11739));
NOR2XL inst_cellmath__62_0_I1484 (.Y(N5310), .A(N5207), .B(N5176));
INVXL inst_cellmath__62_0_I1485 (.Y(N5280), .A(N454));
NOR2XL inst_cellmath__62_0_I1486 (.Y(N5251), .A(N5280), .B(N5382));
NOR2XL inst_cellmath__62_0_I1487 (.Y(N5403), .A(N5280), .B(N5117));
NOR2XL inst_cellmath__62_0_I1488 (.Y(N5210), .A(N5280), .B(N5188));
NOR2XL inst_cellmath__62_0_I1489 (.Y(N5360), .A(N5280), .B(N5261));
NOR2XL inst_cellmath__62_0_I1490 (.Y(N5168), .A(N5280), .B(N5336));
NOR2XL inst_cellmath__62_0_I1491 (.Y(N5314), .A(N5280), .B(N5074));
NOR2XL inst_cellmath__62_0_I1492 (.Y(N5124), .A(N5280), .B(N5148));
NOR2XL inst_cellmath__62_0_I1493 (.Y(N5270), .A(N5280), .B(N5221));
NOR2XL inst_cellmath__62_0_I1494 (.Y(N5081), .A(N5280), .B(N5294));
NOR2XL inst_cellmath__62_0_I1495 (.Y(N5231), .A(N5280), .B(N5367));
NOR2XL inst_cellmath__62_0_I1496 (.Y(N5379), .A(N5280), .B(N11739));
NOR2XL inst_cellmath__62_0_I1497 (.Y(N5185), .A(N5280), .B(N5176));
INVXL inst_cellmath__62_0_I1498 (.Y(N5357), .A(N455));
NOR2XL inst_cellmath__62_0_I1499 (.Y(N5131), .A(N5357), .B(N5382));
NOR2XL inst_cellmath__62_0_I1500 (.Y(N5276), .A(N5357), .B(N5117));
NOR2XL inst_cellmath__62_0_I1501 (.Y(N5085), .A(N5357), .B(N5188));
NOR2XL inst_cellmath__62_0_I1502 (.Y(N5233), .A(N5357), .B(N5261));
NOR2XL inst_cellmath__62_0_I1503 (.Y(N5384), .A(N5357), .B(N5336));
NOR2XL inst_cellmath__62_0_I1504 (.Y(N5191), .A(N5357), .B(N5074));
NOR2XL inst_cellmath__62_0_I1505 (.Y(N5339), .A(N5357), .B(N5148));
NOR2XL inst_cellmath__62_0_I1506 (.Y(N5150), .A(N5357), .B(N5221));
NOR2XL inst_cellmath__62_0_I1507 (.Y(N5297), .A(N5357), .B(N5294));
NOR2XL inst_cellmath__62_0_I1508 (.Y(N5106), .A(N5357), .B(N5367));
NOR2XL inst_cellmath__62_0_I1509 (.Y(N5249), .A(N5357), .B(N11739));
NOR2XL inst_cellmath__62_0_I1510 (.Y(N5401), .A(N5357), .B(N5176));
INVXL inst_cellmath__62_0_I1511 (.Y(N5088), .A(N456));
NOR2XL inst_cellmath__62_0_I1512 (.Y(N5344), .A(N5088), .B(N5382));
NOR2XL inst_cellmath__62_0_I1513 (.Y(N5156), .A(N5088), .B(N5117));
NOR2XL inst_cellmath__62_0_I1514 (.Y(N5301), .A(N5088), .B(N5188));
NOR2XL inst_cellmath__62_0_I1515 (.Y(N5110), .A(N5088), .B(N5261));
NOR2XL inst_cellmath__62_0_I1516 (.Y(N5256), .A(N5088), .B(N5336));
NOR2XL inst_cellmath__62_0_I1517 (.Y(N5068), .A(N5088), .B(N5074));
NOR2XL inst_cellmath__62_0_I1518 (.Y(N5214), .A(N5088), .B(N5148));
NOR2XL inst_cellmath__62_0_I1519 (.Y(N5363), .A(N5088), .B(N5221));
NOR2XL inst_cellmath__62_0_I1520 (.Y(N5173), .A(N5088), .B(N5294));
NOR2XL inst_cellmath__62_0_I1521 (.Y(N5318), .A(N5088), .B(N5367));
NOR2XL inst_cellmath__62_0_I1522 (.Y(N5127), .A(N5088), .B(N11739));
NOR2XL inst_cellmath__62_0_I1523 (.Y(N5274), .A(N5088), .B(N5176));
INVXL inst_cellmath__62_0_I1524 (.Y(N5166), .A(N457));
NOR2XL inst_cellmath__62_0_I1525 (.Y(N5222), .A(N5166), .B(N5382));
NOR2XL inst_cellmath__62_0_I1526 (.Y(N5368), .A(N5166), .B(N5117));
NOR2XL inst_cellmath__62_0_I1527 (.Y(N5177), .A(N5166), .B(N5188));
NOR2XL inst_cellmath__62_0_I1528 (.Y(N5325), .A(N5166), .B(N5261));
NOR2XL inst_cellmath__62_0_I1529 (.Y(N5135), .A(N5166), .B(N5336));
NOR2XL inst_cellmath__62_0_I1530 (.Y(N5281), .A(N5166), .B(N5074));
NOR2XL inst_cellmath__62_0_I1531 (.Y(N5089), .A(N5166), .B(N5148));
NOR2XL inst_cellmath__62_0_I1532 (.Y(N5237), .A(N5166), .B(N5221));
NOR2XL inst_cellmath__62_0_I1533 (.Y(N5387), .A(N5166), .B(N5294));
NOR2XL inst_cellmath__62_0_I1534 (.Y(N5195), .A(N5166), .B(N5367));
NOR2XL inst_cellmath__62_0_I1535 (.Y(N5341), .A(N5166), .B(N11739));
NOR2XL inst_cellmath__62_0_I1536 (.Y(N5154), .A(N5166), .B(N5176));
OR2XL inst_cellmath__62_0_I5063 (.Y(N5236), .A(a_man[22]), .B(N3467));
NOR2XL inst_cellmath__62_0_I1538 (.Y(N5096), .A(N5236), .B(N5382));
NOR2XL inst_cellmath__62_0_I1539 (.Y(N5242), .A(N5236), .B(N5117));
NOR2XL inst_cellmath__62_0_I1540 (.Y(N5391), .A(N5236), .B(N5188));
NOR2XL inst_cellmath__62_0_I1541 (.Y(N5200), .A(N5236), .B(N5261));
NOR2XL inst_cellmath__62_0_I1542 (.Y(N5347), .A(N5236), .B(N5336));
NOR2XL inst_cellmath__62_0_I1543 (.Y(N5159), .A(N5236), .B(N5074));
NOR2XL inst_cellmath__62_0_I1544 (.Y(N5305), .A(N5236), .B(N5148));
NOR2XL inst_cellmath__62_0_I1545 (.Y(N5115), .A(N5236), .B(N5221));
NOR2XL inst_cellmath__62_0_I1546 (.Y(N5260), .A(N5236), .B(N5294));
NOR2XL inst_cellmath__62_0_I1547 (.Y(N5072), .A(N5236), .B(N5367));
NOR2XL inst_cellmath__62_0_I1548 (.Y(N5219), .A(N5236), .B(N11739));
NOR2XL inst_cellmath__62_0_I1549 (.Y(inst_cellmath__62__W0[24]), .A(N5236), .B(N5176));
ADDHX1 inst_cellmath__62_0_I1550 (.CO(N5323), .S(inst_cellmath__62__W1[6]), .A(N5289), .B(N5158));
ADDHX1 inst_cellmath__62_0_I1551 (.CO(N5133), .S(inst_cellmath__62__W0[7]), .A(N5165), .B(N5302));
ADDFX1 inst_cellmath__62_0_I1552 (.CO(N5279), .S(inst_cellmath__62__W1[7]), .A(N5369), .B(N5097), .CI(N5323));
ADDHX1 inst_cellmath__62_0_I1553 (.CO(N5087), .S(N5356), .A(N5381), .B(N5178));
ADDFX1 inst_cellmath__62_0_I1554 (.CO(N5235), .S(inst_cellmath__62__W0[8]), .A(N5112), .B(N5311), .CI(N5243));
ADDFX1 inst_cellmath__62_0_I1555 (.CO(inst_cellmath__62__W0[9]), .S(inst_cellmath__62__W1[8]), .A(N5356), .B(N5133), .CI(N5279));
ADDHX1 inst_cellmath__62_0_I1556 (.CO(N5194), .S(N5121), .A(N5251), .B(N5393));
ADDFX1 inst_cellmath__62_0_I1557 (.CO(N5340), .S(N5266), .A(N5258), .B(N5187), .CI(N5122));
ADDFX1 inst_cellmath__62_0_I1558 (.CO(N5153), .S(N5077), .A(N5087), .B(N5327), .CI(N5121));
ADDFX1 inst_cellmath__62_0_I1559 (.CO(inst_cellmath__62__W0[10]), .S(inst_cellmath__62__W1[9]), .A(N5266), .B(N5235), .CI(N5077));
ADDHX1 inst_cellmath__62_0_I1560 (.CO(N5108), .S(N5373), .A(N5131), .B(N5267));
ADDFX1 inst_cellmath__62_0_I1561 (.CO(N5252), .S(N5180), .A(N5136), .B(N5403), .CI(N5335));
ADDFX1 inst_cellmath__62_0_I1562 (.CO(N5064), .S(N5329), .A(N5069), .B(N5201), .CI(N5194));
ADDFX1 inst_cellmath__62_0_I1563 (.CO(N5211), .S(N5140), .A(N5340), .B(N5373), .CI(N5180));
ADDFX1 inst_cellmath__62_0_I1564 (.CO(inst_cellmath__62__W0[11]), .S(inst_cellmath__62__W1[10]), .A(N5329), .B(N5153), .CI(N5140));
ADDHX1 inst_cellmath__62_0_I1565 (.CO(N5169), .S(N5093), .A(N5344), .B(N5147));
ADDFX1 inst_cellmath__62_0_I1566 (.CO(N5315), .S(N5240), .A(N5348), .B(N5276), .CI(N5210));
ADDFX1 inst_cellmath__62_0_I1567 (.CO(N5125), .S(N5390), .A(N5282), .B(N5078), .CI(N5216));
ADDFX1 inst_cellmath__62_0_I1568 (.CO(N5271), .S(N5199), .A(N5093), .B(N5108), .CI(N5252));
ADDFX1 inst_cellmath__62_0_I1569 (.CO(N5082), .S(N5346), .A(N5240), .B(N5064), .CI(N5390));
ADDFX1 inst_cellmath__62_0_I1570 (.CO(inst_cellmath__62__W0[12]), .S(inst_cellmath__62__W1[11]), .A(N5211), .B(N5199), .CI(N5346));
ADDHX1 inst_cellmath__62_0_I1571 (.CO(N5380), .S(N5304), .A(N5222), .B(N5360));
ADDFX1 inst_cellmath__62_0_I1572 (.CO(N5186), .S(N5114), .A(N5226), .B(N5156), .CI(N5085));
ADDFX1 inst_cellmath__62_0_I1573 (.CO(N5334), .S(N5259), .A(N5160), .B(N5293), .CI(N5365));
ADDFX1 inst_cellmath__62_0_I1574 (.CO(N5146), .S(N5071), .A(N5169), .B(N5091), .CI(N5304));
ADDFX1 inst_cellmath__62_0_I1575 (.CO(N5292), .S(N5218), .A(N5125), .B(N5315), .CI(N5114));
ADDFX1 inst_cellmath__62_0_I1576 (.CO(N5100), .S(N5366), .A(N5259), .B(N5271), .CI(N5071));
ADDFX1 inst_cellmath__62_0_I1577 (.CO(inst_cellmath__62__W0[13]), .S(inst_cellmath__62__W1[12]), .A(N5218), .B(N5082), .CI(N5366));
ADDHX1 inst_cellmath__62_0_I1578 (.CO(N5397), .S(N5322), .A(N5096), .B(N5233));
ADDFX1 inst_cellmath__62_0_I1579 (.CO(N5205), .S(N5132), .A(N5101), .B(N5368), .CI(N5301));
ADDFX1 inst_cellmath__62_0_I1580 (.CO(N5354), .S(N5278), .A(N5374), .B(N5168), .CI(N5238));
ADDFX1 inst_cellmath__62_0_I1581 (.CO(N5163), .S(N5086), .A(N5380), .B(N5306), .CI(N5174));
ADDFX1 inst_cellmath__62_0_I1582 (.CO(N5309), .S(N5234), .A(N5186), .B(N5322), .CI(N5334));
ADDFX1 inst_cellmath__62_0_I1583 (.CO(N5120), .S(N5386), .A(N5146), .B(N5132), .CI(N5278));
ADDFX1 inst_cellmath__62_0_I1584 (.CO(N5265), .S(N5192), .A(N5292), .B(N5086), .CI(N5234));
ADDFX1 inst_cellmath__62_0_I1585 (.CO(inst_cellmath__62__W0[14]), .S(inst_cellmath__62__W1[13]), .A(N5386), .B(N5100), .CI(N5192));
ADDFX1 inst_cellmath__62_0_I1586 (.CO(N5225), .S(N5152), .A(N5314), .B(N5242), .CI(N5177));
ADDFX1 inst_cellmath__62_0_I1587 (.CO(N5372), .S(N5298), .A(N5110), .B(N5384), .CI(N5247));
ADDFX1 inst_cellmath__62_0_I1588 (.CO(N5179), .S(N5107), .A(N5388), .B(N5116), .CI(N5181));
ADDFX1 inst_cellmath__62_0_I1589 (.CO(N5328), .S(N5250), .A(N5320), .B(N5397), .CI(N5205));
ADDFX1 inst_cellmath__62_0_I1590 (.CO(N5139), .S(N5402), .A(N5163), .B(N5354), .CI(N5152));
ADDFX1 inst_cellmath__62_0_I1591 (.CO(N5285), .S(N5209), .A(N5107), .B(N5298), .CI(N5309));
ADDFXL inst_cellmath__62_0_I1592 (.CO(N5092), .S(N5359), .A(N5120), .B(N5250), .CI(N5402));
ADDFX1 inst_cellmath__62_0_I1593 (.CO(inst_cellmath__62__W0[15]), .S(inst_cellmath__62__W1[14]), .A(N5265), .B(N5209), .CI(N5359));
ADDFX1 inst_cellmath__62_0_I1594 (.CO(N5389), .S(N5313), .A(N5256), .B(N5191), .CI(N5325));
ADDFX1 inst_cellmath__62_0_I1595 (.CO(N5198), .S(N5123), .A(N5124), .B(N5391), .CI(N5330));
ADDFX1 inst_cellmath__62_0_I1596 (.CO(N5345), .S(N5269), .A(N5398), .B(N5262), .CI(N5197));
ADDFX1 inst_cellmath__62_0_I1597 (.CO(N5157), .S(N5080), .A(N5225), .B(N5129), .CI(N5372));
ADDFXL inst_cellmath__62_0_I1598 (.CO(N5303), .S(N5230), .A(N5313), .B(N5179), .CI(N5328));
ADDFX1 inst_cellmath__62_0_I1599 (.CO(N5113), .S(N5378), .A(N5269), .B(N5123), .CI(N5139));
ADDFXL inst_cellmath__62_0_I1600 (.CO(N5257), .S(N5184), .A(N5285), .B(N5080), .CI(N5230));
ADDFX1 inst_cellmath__62_0_I1601 (.CO(inst_cellmath__62__W0[16]), .S(inst_cellmath__62__W1[15]), .A(N5378), .B(N5092), .CI(N5184));
ADDHX1 inst_cellmath__62_0_I1602 (.CO(N5217), .S(N5145), .A(N5068), .B(N5339));
ADDFX1 inst_cellmath__62_0_I1603 (.CO(N5364), .S(N5291), .A(N5200), .B(N5135), .CI(N5206));
ADDFX1 inst_cellmath__62_0_I1604 (.CO(N5175), .S(N5099), .A(N5270), .B(N5141), .CI(N5073));
ADDFX1 inst_cellmath__62_0_I1605 (.CO(N5321), .S(N5246), .A(N5145), .B(N5342), .CI(N5389));
ADDFX1 inst_cellmath__62_0_I1606 (.CO(N5128), .S(N5395), .A(N5345), .B(N5198), .CI(N5291));
ADDFX1 inst_cellmath__62_0_I1607 (.CO(N5275), .S(N5203), .A(N5099), .B(N5157), .CI(N5246));
ADDFXL inst_cellmath__62_0_I1608 (.CO(N5083), .S(N5351), .A(N5303), .B(N5113), .CI(N5395));
ADDFHXL inst_cellmath__62_0_I1609 (.CO(inst_cellmath__62__W0[17]), .S(inst_cellmath__62__W1[16]), .A(N5257), .B(N5203), .CI(N5351));
ADDFX1 inst_cellmath__62_0_I1610 (.CO(N5383), .S(N5307), .A(N5347), .B(N5281), .CI(N5214));
ADDFX1 inst_cellmath__62_0_I1611 (.CO(N5189), .S(N5118), .A(N5355), .B(N5081), .CI(N5150));
ADDFX1 inst_cellmath__62_0_I1612 (.CO(N5337), .S(N5263), .A(N5220), .B(N5217), .CI(N5286));
ADDFX1 inst_cellmath__62_0_I1613 (.CO(N5149), .S(N5075), .A(N5175), .B(N5364), .CI(N5307));
ADDFXL inst_cellmath__62_0_I1614 (.CO(N5295), .S(N5223), .A(N5321), .B(N5118), .CI(N5263));
ADDFXL inst_cellmath__62_0_I1615 (.CO(N5104), .S(N5370), .A(N5075), .B(N5128), .CI(N5275));
ADDFX1 inst_cellmath__62_0_I1616 (.CO(inst_cellmath__62__W0[18]), .S(inst_cellmath__62__W1[17]), .A(N5083), .B(N5223), .CI(N5370));
ADDFX1 inst_cellmath__62_0_I1617 (.CO(N5400), .S(N5326), .A(N5089), .B(N5159), .CI(N5297));
ADDFX1 inst_cellmath__62_0_I1618 (.CO(N5208), .S(N5137), .A(N5363), .B(N5231), .CI(N5164));
ADDFX1 inst_cellmath__62_0_I1619 (.CO(N5358), .S(N5283), .A(N5383), .B(N5094), .CI(N5189));
ADDFX1 inst_cellmath__62_0_I1620 (.CO(N5167), .S(N5090), .A(N5326), .B(N5337), .CI(N5137));
ADDFXL inst_cellmath__62_0_I1621 (.CO(N5312), .S(N5239), .A(N5283), .B(N5149), .CI(N5295));
ADDFXL inst_cellmath__62_0_I1622 (.CO(inst_cellmath__62__W0[19]), .S(inst_cellmath__62__W1[18]), .A(N5104), .B(N5090), .CI(N5239));
ADDFX1 inst_cellmath__62_0_I1623 (.CO(N5268), .S(N5196), .A(N5173), .B(N5305), .CI(N5237));
ADDFX1 inst_cellmath__62_0_I1624 (.CO(N5079), .S(N5343), .A(N5379), .B(N5106), .CI(N5310));
ADDFX1 inst_cellmath__62_0_I1625 (.CO(N5228), .S(N5155), .A(N5208), .B(N5400), .CI(N5196));
ADDFX1 inst_cellmath__62_0_I1626 (.CO(N5376), .S(N5299), .A(N5358), .B(N5343), .CI(N5167));
ADDFX1 inst_cellmath__62_0_I1627 (.CO(inst_cellmath__62__W0[20]), .S(inst_cellmath__62__W1[19]), .A(N5312), .B(N5155), .CI(N5299));
ADDFX1 inst_cellmath__62_0_I1628 (.CO(N5332), .S(N5254), .A(N5318), .B(N5387), .CI(N5115));
ADDFX1 inst_cellmath__62_0_I1629 (.CO(N5143), .S(N5066), .A(N5185), .B(N5249), .CI(N5268));
ADDFX1 inst_cellmath__62_0_I1630 (.CO(N5288), .S(N5213), .A(N5254), .B(N5079), .CI(N5066));
ADDFX1 inst_cellmath__62_0_I1631 (.CO(inst_cellmath__62__W0[21]), .S(inst_cellmath__62__W1[20]), .A(N5376), .B(N5228), .CI(N5213));
ADDFX1 inst_cellmath__62_0_I1632 (.CO(N5244), .S(N5171), .A(N5195), .B(N5260), .CI(N5127));
ADDFX1 inst_cellmath__62_0_I1633 (.CO(N5392), .S(N5317), .A(N5332), .B(N5401), .CI(N5171));
ADDFX1 inst_cellmath__62_0_I1634 (.CO(inst_cellmath__62__W1[22]), .S(inst_cellmath__62__W1[21]), .A(N5317), .B(N5143), .CI(N5288));
ADDFX1 inst_cellmath__62_0_I1635 (.CO(N5349), .S(N5272), .A(N5341), .B(N5072), .CI(N5274));
ADDFX1 inst_cellmath__62_0_I1636 (.CO(inst_cellmath__62__W1[23]), .S(inst_cellmath__62__W0[22]), .A(N5272), .B(N5244), .CI(N5392));
ADDFX1 inst_cellmath__62_0_I1637 (.CO(inst_cellmath__62__W1[24]), .S(inst_cellmath__62__W0[23]), .A(N5154), .B(N5219), .CI(N5349));
INVXL inst_cellmath__63_0_I1638 (.Y(N6077), .A(inst_cellmath__51[0]));
INVXL inst_cellmath__63_0_I1639 (.Y(N6533), .A(inst_cellmath__51[1]));
INVXL inst_cellmath__63_0_I1640 (.Y(N6122), .A(inst_cellmath__51[2]));
INVXL inst_cellmath__63_0_I1641 (.Y(N6578), .A(inst_cellmath__51[3]));
INVXL inst_cellmath__63_0_I1642 (.Y(N6168), .A(inst_cellmath__51[4]));
INVXL inst_cellmath__63_0_I1643 (.Y(N5761), .A(inst_cellmath__51[5]));
INVXL inst_cellmath__63_0_I1644 (.Y(N6217), .A(inst_cellmath__51[6]));
INVXL inst_cellmath__63_0_I1645 (.Y(N5810), .A(inst_cellmath__51[7]));
INVXL inst_cellmath__63_0_I1646 (.Y(N6260), .A(inst_cellmath__51[8]));
INVXL inst_cellmath__63_0_I1647 (.Y(N5852), .A(inst_cellmath__51[9]));
INVXL inst_cellmath__63_0_I1648 (.Y(N6305), .A(inst_cellmath__51[10]));
INVXL inst_cellmath__63_0_I1649 (.Y(N5897), .A(inst_cellmath__51[11]));
INVXL inst_cellmath__63_0_I1650 (.Y(N6356), .A(inst_cellmath__51[12]));
INVXL inst_cellmath__63_0_I1651 (.Y(N5947), .A(inst_cellmath__51[13]));
INVXL inst_cellmath__63_0_I1652 (.Y(N6403), .A(inst_cellmath__51[14]));
INVXL inst_cellmath__63_0_I1653 (.Y(N5992), .A(inst_cellmath__51[15]));
INVXL inst_cellmath__63_0_I1654 (.Y(N6446), .A(inst_cellmath__51[16]));
INVXL inst_cellmath__63_0_I1655 (.Y(N6035), .A(inst_cellmath__51[17]));
INVXL inst_cellmath__63_0_I1656 (.Y(N6301), .A(a_man[0]));
NOR2XL inst_cellmath__63_0_I1659 (.Y(N5971), .A(N6301), .B(N6122));
NOR2XL inst_cellmath__63_0_I1660 (.Y(N6349), .A(N6301), .B(N6578));
NOR2XL inst_cellmath__63_0_I1661 (.Y(N5861), .A(N6301), .B(N6168));
NOR2XL inst_cellmath__63_0_I1662 (.Y(N6234), .A(N6301), .B(N5761));
NOR2XL inst_cellmath__63_0_I1663 (.Y(N5750), .A(N6301), .B(N6217));
NOR2XL inst_cellmath__63_0_I1664 (.Y(N6128), .A(N6301), .B(N5810));
NOR2XL inst_cellmath__63_0_I1665 (.Y(N6503), .A(N6301), .B(N6260));
NOR2XL inst_cellmath__63_0_I1666 (.Y(N6018), .A(N6301), .B(N5852));
NOR2XL inst_cellmath__63_0_I1667 (.Y(N6398), .A(N6301), .B(N6305));
NOR2XL inst_cellmath__63_0_I1668 (.Y(N5906), .A(N6301), .B(N5897));
NOR2XL inst_cellmath__63_0_I1669 (.Y(N6282), .A(N6301), .B(N6356));
NOR2XL inst_cellmath__63_0_I1670 (.Y(N5799), .A(N6301), .B(N5947));
NOR2XL inst_cellmath__63_0_I1671 (.Y(N6172), .A(N6301), .B(N6403));
NOR2XL inst_cellmath__63_0_I1672 (.Y(N6550), .A(N6301), .B(N5992));
NOR2XL inst_cellmath__63_0_I1673 (.Y(N6062), .A(N6301), .B(N6446));
NOR2XL inst_cellmath__63_0_I1674 (.Y(N6438), .A(N6301), .B(N6035));
INVXL inst_cellmath__63_0_I1675 (.Y(N6570), .A(a_man[1]));
NOR2XL inst_cellmath__63_0_I1677 (.Y(inst_cellmath__63__W0[2]), .A(N6570), .B(N6533));
NOR2XL inst_cellmath__63_0_I1678 (.Y(N6379), .A(N6570), .B(N6122));
NOR2XL inst_cellmath__63_0_I1679 (.Y(N5889), .A(N6570), .B(N6578));
NOR2XL inst_cellmath__63_0_I1680 (.Y(N6265), .A(N6570), .B(N6168));
NOR2XL inst_cellmath__63_0_I1681 (.Y(N5781), .A(N6570), .B(N5761));
NOR2XL inst_cellmath__63_0_I1682 (.Y(N6154), .A(N6570), .B(N6217));
NOR2XL inst_cellmath__63_0_I1683 (.Y(N6535), .A(N6570), .B(N5810));
NOR2XL inst_cellmath__63_0_I1684 (.Y(N6042), .A(N6570), .B(N6260));
NOR2XL inst_cellmath__63_0_I1685 (.Y(N6422), .A(N6570), .B(N5852));
NOR2XL inst_cellmath__63_0_I1686 (.Y(N5935), .A(N6570), .B(N6305));
NOR2XL inst_cellmath__63_0_I1687 (.Y(N6311), .A(N6570), .B(N5897));
NOR2XL inst_cellmath__63_0_I1688 (.Y(N5826), .A(N6570), .B(N6356));
NOR2XL inst_cellmath__63_0_I1689 (.Y(N6201), .A(N6570), .B(N5947));
NOR2XL inst_cellmath__63_0_I1690 (.Y(N6580), .A(N6570), .B(N6403));
NOR2XL inst_cellmath__63_0_I1691 (.Y(N6088), .A(N6570), .B(N5992));
NOR2XL inst_cellmath__63_0_I1692 (.Y(N6469), .A(N6570), .B(N6446));
NOR2XL inst_cellmath__63_0_I1693 (.Y(N5982), .A(N6570), .B(N6035));
INVXL inst_cellmath__63_0_I1694 (.Y(N5975), .A(a_man[2]));
NOR2XL inst_cellmath__63_0_I1695 (.Y(N6029), .A(N5975), .B(N6077));
NOR2XL inst_cellmath__63_0_I1696 (.Y(N6408), .A(N5975), .B(N6533));
NOR2XL inst_cellmath__63_0_I1697 (.Y(N5918), .A(N5975), .B(N6122));
NOR2XL inst_cellmath__63_0_I1698 (.Y(N6293), .A(N5975), .B(N6578));
NOR2XL inst_cellmath__63_0_I1699 (.Y(N5811), .A(N5975), .B(N6168));
NOR2XL inst_cellmath__63_0_I1700 (.Y(N6186), .A(N5975), .B(N5761));
NOR2XL inst_cellmath__63_0_I1701 (.Y(N6560), .A(N5975), .B(N6217));
NOR2XL inst_cellmath__63_0_I1702 (.Y(N6073), .A(N5975), .B(N5810));
NOR2XL inst_cellmath__63_0_I1703 (.Y(N6452), .A(N5975), .B(N6260));
NOR2XL inst_cellmath__63_0_I1704 (.Y(N5964), .A(N5975), .B(N5852));
NOR2XL inst_cellmath__63_0_I1705 (.Y(N6341), .A(N5975), .B(N6305));
NOR2XL inst_cellmath__63_0_I1706 (.Y(N5853), .A(N5975), .B(N5897));
NOR2XL inst_cellmath__63_0_I1707 (.Y(N6227), .A(N5975), .B(N6356));
NOR2XL inst_cellmath__63_0_I1708 (.Y(N5743), .A(N5975), .B(N5947));
NOR2XL inst_cellmath__63_0_I1709 (.Y(N6118), .A(N5975), .B(N6403));
NOR2XL inst_cellmath__63_0_I1710 (.Y(N6494), .A(N5975), .B(N5992));
NOR2XL inst_cellmath__63_0_I1711 (.Y(N6009), .A(N5975), .B(N6446));
NOR2XL inst_cellmath__63_0_I1712 (.Y(N6389), .A(N5975), .B(N6035));
NOR2XL inst_cellmath__63_0_I1714 (.Y(N6432), .A(N2876), .B(N6077));
NOR2XL inst_cellmath__63_0_I1715 (.Y(N5949), .A(N2876), .B(N6533));
NOR2XL inst_cellmath__63_0_I1716 (.Y(N6325), .A(N2876), .B(N6122));
NOR2XL inst_cellmath__63_0_I1717 (.Y(N5838), .A(N2876), .B(N6578));
NOR2XL inst_cellmath__63_0_I1718 (.Y(N6213), .A(N2876), .B(N6168));
NOR2XL inst_cellmath__63_0_I1719 (.Y(N5730), .A(N2876), .B(N5761));
NOR2XL inst_cellmath__63_0_I1720 (.Y(N6100), .A(N2876), .B(N6217));
NOR2XL inst_cellmath__63_0_I1721 (.Y(N6481), .A(N2876), .B(N5810));
NOR2XL inst_cellmath__63_0_I1722 (.Y(N5994), .A(N2876), .B(N6260));
NOR2XL inst_cellmath__63_0_I1723 (.Y(N6369), .A(N2876), .B(N5852));
NOR2XL inst_cellmath__63_0_I1724 (.Y(N5881), .A(N2876), .B(N6305));
NOR2XL inst_cellmath__63_0_I1725 (.Y(N6256), .A(N2876), .B(N5897));
NOR2XL inst_cellmath__63_0_I1726 (.Y(N5771), .A(N2876), .B(N6356));
NOR2XL inst_cellmath__63_0_I1727 (.Y(N6146), .A(N2876), .B(N5947));
NOR2XL inst_cellmath__63_0_I1728 (.Y(N6525), .A(N2876), .B(N6403));
NOR2XL inst_cellmath__63_0_I1729 (.Y(N6034), .A(N2876), .B(N5992));
NOR2XL inst_cellmath__63_0_I1730 (.Y(N6414), .A(N2876), .B(N6446));
NOR2XL inst_cellmath__63_0_I1731 (.Y(N5929), .A(N2876), .B(N6035));
NOR2XL inst_cellmath__63_0_I1733 (.Y(N5977), .A(N11660), .B(N6077));
NOR2XL inst_cellmath__63_0_I1734 (.Y(N6353), .A(N11660), .B(N6533));
NOR2XL inst_cellmath__63_0_I1735 (.Y(N5865), .A(N11660), .B(N6122));
NOR2XL inst_cellmath__63_0_I1736 (.Y(N6240), .A(N11660), .B(N6578));
NOR2XL inst_cellmath__63_0_I1737 (.Y(N5754), .A(N11660), .B(N6168));
NOR2XL inst_cellmath__63_0_I1738 (.Y(N6132), .A(N11660), .B(N5761));
NOR2XL inst_cellmath__63_0_I1739 (.Y(N6509), .A(N11660), .B(N6217));
NOR2XL inst_cellmath__63_0_I1740 (.Y(N6022), .A(N11661), .B(N5810));
NOR2XL inst_cellmath__63_0_I1741 (.Y(N6400), .A(N11661), .B(N6260));
NOR2XL inst_cellmath__63_0_I1742 (.Y(N5912), .A(N11661), .B(N5852));
NOR2XL inst_cellmath__63_0_I1743 (.Y(N6285), .A(N11661), .B(N6305));
NOR2XL inst_cellmath__63_0_I1744 (.Y(N5802), .A(N11661), .B(N5897));
NOR2XL inst_cellmath__63_0_I1745 (.Y(N6177), .A(N11661), .B(N6356));
NOR2XL inst_cellmath__63_0_I1746 (.Y(N6553), .A(N11661), .B(N5947));
NOR2XL inst_cellmath__63_0_I1747 (.Y(N6065), .A(N11661), .B(N6403));
NOR2XL inst_cellmath__63_0_I1748 (.Y(N6442), .A(N11660), .B(N5992));
NOR2XL inst_cellmath__63_0_I1749 (.Y(N5956), .A(N11660), .B(N6446));
NOR2XL inst_cellmath__63_0_I1750 (.Y(N6333), .A(N11660), .B(N6035));
NOR2XL inst_cellmath__63_0_I1752 (.Y(N6383), .A(N11669), .B(N6077));
NOR2XL inst_cellmath__63_0_I1753 (.Y(N5892), .A(N11669), .B(N6533));
NOR2XL inst_cellmath__63_0_I1754 (.Y(N6268), .A(N11669), .B(N6122));
NOR2XL inst_cellmath__63_0_I1755 (.Y(N5785), .A(N11669), .B(N6578));
NOR2XL inst_cellmath__63_0_I1756 (.Y(N6157), .A(N11669), .B(N6168));
NOR2XL inst_cellmath__63_0_I1757 (.Y(N6538), .A(N11669), .B(N5761));
NOR2XL inst_cellmath__63_0_I1758 (.Y(N6047), .A(N11669), .B(N6217));
NOR2XL inst_cellmath__63_0_I1759 (.Y(N6424), .A(N11669), .B(N5810));
NOR2XL inst_cellmath__63_0_I1760 (.Y(N5939), .A(N11669), .B(N6260));
NOR2XL inst_cellmath__63_0_I1761 (.Y(N6316), .A(N11669), .B(N5852));
NOR2XL inst_cellmath__63_0_I1762 (.Y(N5830), .A(N11669), .B(N6305));
NOR2XL inst_cellmath__63_0_I1763 (.Y(N6205), .A(N11669), .B(N5897));
NOR2XL inst_cellmath__63_0_I1764 (.Y(N5724), .A(N11669), .B(N6356));
NOR2XL inst_cellmath__63_0_I1765 (.Y(N6092), .A(N11669), .B(N5947));
NOR2XL inst_cellmath__63_0_I1766 (.Y(N6473), .A(N11669), .B(N6403));
NOR2XL inst_cellmath__63_0_I1767 (.Y(N5985), .A(N11669), .B(N5992));
NOR2XL inst_cellmath__63_0_I1768 (.Y(N6361), .A(N11669), .B(N6446));
NOR2XL inst_cellmath__63_0_I1769 (.Y(N5873), .A(N11669), .B(N6035));
NOR2XL inst_cellmath__63_0_I1771 (.Y(N5921), .A(N2773), .B(N6077));
NOR2XL inst_cellmath__63_0_I1772 (.Y(N6295), .A(N2773), .B(N6533));
NOR2XL inst_cellmath__63_0_I1773 (.Y(N5813), .A(N2773), .B(N6122));
NOR2XL inst_cellmath__63_0_I1774 (.Y(N6189), .A(N2773), .B(N6578));
NOR2XL inst_cellmath__63_0_I1775 (.Y(N6562), .A(N2773), .B(N6168));
NOR2XL inst_cellmath__63_0_I1776 (.Y(N6076), .A(N2773), .B(N5761));
NOR2XL inst_cellmath__63_0_I1777 (.Y(N6455), .A(N2773), .B(N6217));
NOR2XL inst_cellmath__63_0_I1778 (.Y(N5966), .A(N2773), .B(N5810));
NOR2XL inst_cellmath__63_0_I1779 (.Y(N6344), .A(N2773), .B(N6260));
NOR2XL inst_cellmath__63_0_I1780 (.Y(N5856), .A(N2773), .B(N5852));
NOR2XL inst_cellmath__63_0_I1781 (.Y(N6229), .A(N2773), .B(N6305));
NOR2XL inst_cellmath__63_0_I1782 (.Y(N5745), .A(N2773), .B(N5897));
NOR2XL inst_cellmath__63_0_I1783 (.Y(N6121), .A(N2773), .B(N6356));
NOR2XL inst_cellmath__63_0_I1784 (.Y(N6497), .A(N2773), .B(N5947));
NOR2XL inst_cellmath__63_0_I1785 (.Y(N6012), .A(N2773), .B(N6403));
NOR2XL inst_cellmath__63_0_I1786 (.Y(N6392), .A(N2773), .B(N5992));
NOR2XL inst_cellmath__63_0_I1787 (.Y(N5900), .A(N2773), .B(N6446));
NOR2XL inst_cellmath__63_0_I1788 (.Y(N6276), .A(N2773), .B(N6035));
NOR2XL inst_cellmath__63_0_I1790 (.Y(N6328), .A(N11688), .B(N6077));
NOR2XL inst_cellmath__63_0_I1791 (.Y(N5841), .A(N11688), .B(N6533));
NOR2XL inst_cellmath__63_0_I1792 (.Y(N6216), .A(N11688), .B(N6122));
NOR2XL inst_cellmath__63_0_I1793 (.Y(N5733), .A(N11688), .B(N6578));
NOR2XL inst_cellmath__63_0_I1794 (.Y(N6103), .A(N11688), .B(N6168));
NOR2XL inst_cellmath__63_0_I1795 (.Y(N6484), .A(N11688), .B(N5761));
NOR2XL inst_cellmath__63_0_I1796 (.Y(N5997), .A(N11688), .B(N6217));
NOR2XL inst_cellmath__63_0_I1797 (.Y(N6373), .A(N11688), .B(N5810));
NOR2XL inst_cellmath__63_0_I1798 (.Y(N5883), .A(N11688), .B(N6260));
NOR2XL inst_cellmath__63_0_I1799 (.Y(N6259), .A(N11688), .B(N5852));
NOR2XL inst_cellmath__63_0_I1800 (.Y(N5775), .A(N11688), .B(N6305));
NOR2XL inst_cellmath__63_0_I1801 (.Y(N6148), .A(N11688), .B(N5897));
NOR2XL inst_cellmath__63_0_I1802 (.Y(N6528), .A(N11688), .B(N6356));
NOR2XL inst_cellmath__63_0_I1803 (.Y(N6038), .A(N11688), .B(N5947));
NOR2XL inst_cellmath__63_0_I1804 (.Y(N6416), .A(N11688), .B(N6403));
NOR2XL inst_cellmath__63_0_I1805 (.Y(N5930), .A(N11688), .B(N5992));
NOR2XL inst_cellmath__63_0_I1806 (.Y(N6304), .A(N11688), .B(N6446));
NOR2XL inst_cellmath__63_0_I1807 (.Y(N5820), .A(N11688), .B(N6035));
NOR2XL inst_cellmath__63_0_I1809 (.Y(N5867), .A(N11693), .B(N6077));
NOR2XL inst_cellmath__63_0_I1810 (.Y(N6243), .A(N11693), .B(N6533));
NOR2XL inst_cellmath__63_0_I1811 (.Y(N5756), .A(N11693), .B(N6122));
NOR2XL inst_cellmath__63_0_I1812 (.Y(N6134), .A(N11693), .B(N6578));
NOR2XL inst_cellmath__63_0_I1813 (.Y(N6512), .A(N11693), .B(N6168));
NOR2XL inst_cellmath__63_0_I1814 (.Y(N6024), .A(N11693), .B(N5761));
NOR2XL inst_cellmath__63_0_I1815 (.Y(N6401), .A(N11693), .B(N6217));
NOR2XL inst_cellmath__63_0_I1816 (.Y(N5915), .A(N11693), .B(N5810));
NOR2XL inst_cellmath__63_0_I1817 (.Y(N6287), .A(N11693), .B(N6260));
NOR2XL inst_cellmath__63_0_I1818 (.Y(N5804), .A(N11693), .B(N5852));
NOR2XL inst_cellmath__63_0_I1819 (.Y(N6180), .A(N11693), .B(N6305));
NOR2XL inst_cellmath__63_0_I1820 (.Y(N6555), .A(N11693), .B(N5897));
NOR2XL inst_cellmath__63_0_I1821 (.Y(N6067), .A(N11693), .B(N6356));
NOR2XL inst_cellmath__63_0_I1822 (.Y(N6445), .A(N11693), .B(N5947));
NOR2XL inst_cellmath__63_0_I1823 (.Y(N5958), .A(N11693), .B(N6403));
NOR2XL inst_cellmath__63_0_I1824 (.Y(N6335), .A(N11693), .B(N5992));
NOR2XL inst_cellmath__63_0_I1825 (.Y(N5848), .A(N11697), .B(N6446));
NOR2XL inst_cellmath__63_0_I1826 (.Y(N6223), .A(N11697), .B(N6035));
NOR2XL inst_cellmath__63_0_I1828 (.Y(N6270), .A(N11706), .B(N6077));
NOR2XL inst_cellmath__63_0_I1829 (.Y(N5787), .A(N11706), .B(N6533));
NOR2XL inst_cellmath__63_0_I1830 (.Y(N6158), .A(N11706), .B(N6122));
NOR2XL inst_cellmath__63_0_I1831 (.Y(N6540), .A(N11706), .B(N6578));
NOR2XL inst_cellmath__63_0_I1832 (.Y(N6049), .A(N11706), .B(N6168));
NOR2XL inst_cellmath__63_0_I1833 (.Y(N6425), .A(N11706), .B(N5761));
NOR2XL inst_cellmath__63_0_I1834 (.Y(N5941), .A(N11706), .B(N6217));
NOR2XL inst_cellmath__63_0_I1835 (.Y(N6318), .A(N11706), .B(N5810));
NOR2XL inst_cellmath__63_0_I1836 (.Y(N5831), .A(N11706), .B(N6260));
NOR2XL inst_cellmath__63_0_I1837 (.Y(N6206), .A(N11706), .B(N5852));
NOR2XL inst_cellmath__63_0_I1838 (.Y(N5726), .A(N11706), .B(N6305));
NOR2XL inst_cellmath__63_0_I1839 (.Y(N6093), .A(N11706), .B(N5897));
NOR2XL inst_cellmath__63_0_I1840 (.Y(N6475), .A(N11706), .B(N6356));
NOR2XL inst_cellmath__63_0_I1841 (.Y(N5987), .A(N11706), .B(N5947));
NOR2XL inst_cellmath__63_0_I1842 (.Y(N6363), .A(N11706), .B(N6403));
NOR2XL inst_cellmath__63_0_I1843 (.Y(N5875), .A(N11706), .B(N5992));
NOR2XL inst_cellmath__63_0_I1844 (.Y(N6250), .A(N11706), .B(N6446));
NOR2XL inst_cellmath__63_0_I1845 (.Y(N5765), .A(N11706), .B(N6035));
NOR2XL inst_cellmath__63_0_I1847 (.Y(N5815), .A(N11708), .B(N6077));
NOR2XL inst_cellmath__63_0_I1848 (.Y(N6191), .A(N11708), .B(N6533));
NOR2XL inst_cellmath__63_0_I1849 (.Y(N6564), .A(N11708), .B(N6122));
NOR2XL inst_cellmath__63_0_I1850 (.Y(N6079), .A(N11708), .B(N6578));
NOR2XL inst_cellmath__63_0_I1851 (.Y(N6457), .A(N11708), .B(N6168));
NOR2XL inst_cellmath__63_0_I1852 (.Y(N5968), .A(N11708), .B(N5761));
NOR2XL inst_cellmath__63_0_I1853 (.Y(N6346), .A(N11708), .B(N6217));
NOR2XL inst_cellmath__63_0_I1854 (.Y(N5858), .A(N11708), .B(N5810));
NOR2XL inst_cellmath__63_0_I1855 (.Y(N6232), .A(N11708), .B(N6260));
NOR2XL inst_cellmath__63_0_I1856 (.Y(N5747), .A(N11708), .B(N5852));
NOR2XL inst_cellmath__63_0_I1857 (.Y(N6124), .A(N11708), .B(N6305));
NOR2XL inst_cellmath__63_0_I1858 (.Y(N6501), .A(N11708), .B(N5897));
NOR2XL inst_cellmath__63_0_I1859 (.Y(N6014), .A(N11708), .B(N6356));
NOR2XL inst_cellmath__63_0_I1860 (.Y(N6394), .A(N11708), .B(N5947));
NOR2XL inst_cellmath__63_0_I1861 (.Y(N5904), .A(N11708), .B(N6403));
NOR2XL inst_cellmath__63_0_I1862 (.Y(N6278), .A(N11708), .B(N5992));
NOR2XL inst_cellmath__63_0_I1863 (.Y(N5795), .A(N11708), .B(N6446));
NOR2XL inst_cellmath__63_0_I1864 (.Y(N6170), .A(N11708), .B(N6035));
NOR2XL inst_cellmath__63_0_I1866 (.Y(N6219), .A(N11719), .B(N6077));
NOR2XL inst_cellmath__63_0_I1867 (.Y(N5735), .A(N11719), .B(N6533));
NOR2XL inst_cellmath__63_0_I1868 (.Y(N6106), .A(N11719), .B(N6122));
NOR2XL inst_cellmath__63_0_I1869 (.Y(N6486), .A(N11719), .B(N6578));
NOR2XL inst_cellmath__63_0_I1870 (.Y(N6000), .A(N11719), .B(N6168));
NOR2XL inst_cellmath__63_0_I1871 (.Y(N6376), .A(N11719), .B(N5761));
NOR2XL inst_cellmath__63_0_I1872 (.Y(N5886), .A(N11719), .B(N6217));
NOR2XL inst_cellmath__63_0_I1873 (.Y(N6262), .A(N11719), .B(N5810));
NOR2XL inst_cellmath__63_0_I1874 (.Y(N5778), .A(N11719), .B(N6260));
NOR2XL inst_cellmath__63_0_I1875 (.Y(N6151), .A(N11719), .B(N5852));
NOR2XL inst_cellmath__63_0_I1876 (.Y(N6531), .A(N11719), .B(N6305));
NOR2XL inst_cellmath__63_0_I1877 (.Y(N6039), .A(N11719), .B(N5897));
NOR2XL inst_cellmath__63_0_I1878 (.Y(N6419), .A(N11719), .B(N6356));
NOR2XL inst_cellmath__63_0_I1879 (.Y(N5933), .A(N11719), .B(N5947));
NOR2XL inst_cellmath__63_0_I1880 (.Y(N6308), .A(N11719), .B(N6403));
NOR2XL inst_cellmath__63_0_I1881 (.Y(N5823), .A(N11719), .B(N5992));
NOR2XL inst_cellmath__63_0_I1882 (.Y(N6198), .A(N11719), .B(N6446));
NOR2XL inst_cellmath__63_0_I1883 (.Y(N6576), .A(N11719), .B(N6035));
NOR2XL inst_cellmath__63_0_I1885 (.Y(N5759), .A(N11728), .B(N6077));
NOR2XL inst_cellmath__63_0_I1886 (.Y(N6138), .A(N11728), .B(N6533));
NOR2XL inst_cellmath__63_0_I1887 (.Y(N6515), .A(N11728), .B(N6122));
NOR2XL inst_cellmath__63_0_I1888 (.Y(N6027), .A(N11728), .B(N6578));
NOR2XL inst_cellmath__63_0_I1889 (.Y(N6406), .A(N11728), .B(N6168));
NOR2XL inst_cellmath__63_0_I1890 (.Y(N5916), .A(N11728), .B(N5761));
NOR2XL inst_cellmath__63_0_I1891 (.Y(N6290), .A(N11728), .B(N6217));
NOR2XL inst_cellmath__63_0_I1892 (.Y(N5808), .A(N11728), .B(N5810));
NOR2XL inst_cellmath__63_0_I1893 (.Y(N6183), .A(N11728), .B(N6260));
NOR2XL inst_cellmath__63_0_I1894 (.Y(N6558), .A(N11728), .B(N5852));
NOR2XL inst_cellmath__63_0_I1895 (.Y(N6071), .A(N11728), .B(N6305));
NOR2XL inst_cellmath__63_0_I1896 (.Y(N6449), .A(N11728), .B(N5897));
NOR2XL inst_cellmath__63_0_I1897 (.Y(N5961), .A(N11728), .B(N6356));
NOR2XL inst_cellmath__63_0_I1898 (.Y(N6338), .A(N11728), .B(N5947));
NOR2XL inst_cellmath__63_0_I1899 (.Y(N5850), .A(N11728), .B(N6403));
NOR2XL inst_cellmath__63_0_I1900 (.Y(N6225), .A(N11728), .B(N5992));
NOR2XL inst_cellmath__63_0_I1901 (.Y(N5740), .A(N11728), .B(N6446));
NOR2XL inst_cellmath__63_0_I1902 (.Y(N6116), .A(N11728), .B(N6035));
NOR2XL inst_cellmath__63_0_I1904 (.Y(N6162), .A(N2705), .B(N6077));
NOR2XL inst_cellmath__63_0_I1905 (.Y(N6543), .A(N2705), .B(N6533));
NOR2XL inst_cellmath__63_0_I1906 (.Y(N6052), .A(N2705), .B(N6122));
NOR2XL inst_cellmath__63_0_I1907 (.Y(N6429), .A(N2705), .B(N6578));
NOR2XL inst_cellmath__63_0_I1908 (.Y(N5944), .A(N2705), .B(N6168));
NOR2XL inst_cellmath__63_0_I1909 (.Y(N6321), .A(N2705), .B(N5761));
NOR2XL inst_cellmath__63_0_I1910 (.Y(N5835), .A(N2705), .B(N6217));
NOR2XL inst_cellmath__63_0_I1911 (.Y(N6209), .A(N2705), .B(N5810));
NOR2XL inst_cellmath__63_0_I1912 (.Y(N5728), .A(N2705), .B(N6260));
NOR2XL inst_cellmath__63_0_I1913 (.Y(N6097), .A(N2705), .B(N5852));
NOR2XL inst_cellmath__63_0_I1914 (.Y(N6477), .A(N2705), .B(N6305));
NOR2XL inst_cellmath__63_0_I1915 (.Y(N5989), .A(N2705), .B(N5897));
NOR2XL inst_cellmath__63_0_I1916 (.Y(N6366), .A(N2705), .B(N6356));
NOR2XL inst_cellmath__63_0_I1917 (.Y(N5877), .A(N2705), .B(N5947));
NOR2XL inst_cellmath__63_0_I1918 (.Y(N6252), .A(N2705), .B(N6403));
NOR2XL inst_cellmath__63_0_I1919 (.Y(N5768), .A(N2705), .B(N5992));
NOR2XL inst_cellmath__63_0_I1920 (.Y(N6143), .A(N2705), .B(N6446));
NOR2XL inst_cellmath__63_0_I1921 (.Y(N6522), .A(N2705), .B(N6035));
NOR2XL inst_cellmath__63_0_I1923 (.Y(N6567), .A(N2777), .B(N6077));
NOR2XL inst_cellmath__63_0_I1924 (.Y(N6081), .A(N2777), .B(N6533));
NOR2XL inst_cellmath__63_0_I1925 (.Y(N6459), .A(N2777), .B(N6122));
NOR2XL inst_cellmath__63_0_I1926 (.Y(N5972), .A(N2777), .B(N6578));
NOR2XL inst_cellmath__63_0_I1927 (.Y(N6348), .A(N2777), .B(N6168));
NOR2XL inst_cellmath__63_0_I1928 (.Y(N5860), .A(N2777), .B(N5761));
NOR2XL inst_cellmath__63_0_I1929 (.Y(N6235), .A(N2777), .B(N6217));
NOR2XL inst_cellmath__63_0_I1930 (.Y(N5749), .A(N2777), .B(N5810));
NOR2XL inst_cellmath__63_0_I1931 (.Y(N6127), .A(N2777), .B(N6260));
NOR2XL inst_cellmath__63_0_I1932 (.Y(N6504), .A(N2777), .B(N5852));
NOR2XL inst_cellmath__63_0_I1933 (.Y(N6017), .A(N2777), .B(N6305));
NOR2XL inst_cellmath__63_0_I1934 (.Y(N6397), .A(N2777), .B(N5897));
NOR2XL inst_cellmath__63_0_I1935 (.Y(N5907), .A(N2777), .B(N6356));
NOR2XL inst_cellmath__63_0_I1936 (.Y(N6281), .A(N2777), .B(N5947));
NOR2XL inst_cellmath__63_0_I1937 (.Y(N5798), .A(N2777), .B(N6403));
NOR2XL inst_cellmath__63_0_I1938 (.Y(N6173), .A(N2777), .B(N5992));
NOR2XL inst_cellmath__63_0_I1939 (.Y(N6549), .A(N2777), .B(N6446));
NOR2XL inst_cellmath__63_0_I1940 (.Y(N6061), .A(N2777), .B(N6035));
NAND2XL inst_cellmath__63_0_I1941 (.Y(N6108), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[0]));
NAND2XL inst_cellmath__63_0_I1942 (.Y(N6488), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[1]));
NAND2XL inst_cellmath__63_0_I1943 (.Y(N6002), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[2]));
NAND2XL inst_cellmath__63_0_I1944 (.Y(N6378), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[3]));
NAND2XL inst_cellmath__63_0_I1945 (.Y(N5888), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[4]));
NAND2XL inst_cellmath__63_0_I1946 (.Y(N6264), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[5]));
NAND2XL inst_cellmath__63_0_I1947 (.Y(N5780), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[6]));
NAND2XL inst_cellmath__63_0_I1948 (.Y(N6153), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[7]));
NAND2XL inst_cellmath__63_0_I1949 (.Y(N6534), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[8]));
NAND2XL inst_cellmath__63_0_I1950 (.Y(N6041), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[9]));
NAND2XL inst_cellmath__63_0_I1951 (.Y(N6421), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[10]));
NAND2XL inst_cellmath__63_0_I1952 (.Y(N5934), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[11]));
NAND2XL inst_cellmath__63_0_I1953 (.Y(N6310), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[12]));
NAND2XL inst_cellmath__63_0_I1954 (.Y(N5825), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[13]));
NAND2XL inst_cellmath__63_0_I1955 (.Y(N6200), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[14]));
NAND2XL inst_cellmath__63_0_I1956 (.Y(N6579), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[15]));
NAND2XL inst_cellmath__63_0_I1957 (.Y(N6087), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[16]));
NAND2XL inst_cellmath__63_0_I1958 (.Y(N6468), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[17]));
ADDHX1 inst_cellmath__63_0_I1959 (.CO(N6104), .S(inst_cellmath__63__W1[2]), .A(N5971), .B(N6029));
ADDHX1 inst_cellmath__63_0_I1960 (.CO(N6485), .S(inst_cellmath__63__W0[3]), .A(N6379), .B(N6408));
ADDFX1 inst_cellmath__63_0_I1961 (.CO(N5998), .S(inst_cellmath__63__W1[3]), .A(N6432), .B(N6349), .CI(N6104));
ADDHX1 inst_cellmath__63_0_I1962 (.CO(N6374), .S(N6185), .A(N5918), .B(N5949));
ADDFX1 inst_cellmath__63_0_I1963 (.CO(N5884), .S(inst_cellmath__63__W0[4]), .A(N5861), .B(N5889), .CI(N5977));
ADDFX1 inst_cellmath__63_0_I1964 (.CO(inst_cellmath__63__W0[5]), .S(inst_cellmath__63__W1[4]), .A(N6185), .B(N6485), .CI(N5998));
ADDHX1 inst_cellmath__63_0_I1965 (.CO(N5776), .S(N6451), .A(N6234), .B(N6383));
ADDFX1 inst_cellmath__63_0_I1966 (.CO(N6149), .S(N5963), .A(N6265), .B(N6325), .CI(N6293));
ADDFX1 inst_cellmath__63_0_I1967 (.CO(N6529), .S(N6340), .A(N6374), .B(N6353), .CI(N6451));
ADDFX1 inst_cellmath__63_0_I1968 (.CO(inst_cellmath__63__W0[6]), .S(inst_cellmath__63__W1[5]), .A(N5963), .B(N5884), .CI(N6340));
ADDHX1 inst_cellmath__63_0_I1969 (.CO(N6417), .S(N6228), .A(N5781), .B(N5921));
ADDFX1 inst_cellmath__63_0_I1970 (.CO(N5931), .S(N5742), .A(N5811), .B(N5865), .CI(N5838));
ADDFX1 inst_cellmath__63_0_I1971 (.CO(N6306), .S(N6117), .A(N5892), .B(N5750), .CI(N5776));
ADDFX1 inst_cellmath__63_0_I1972 (.CO(N5821), .S(N6495), .A(N6228), .B(N6149), .CI(N5742));
ADDFX1 inst_cellmath__63_0_I1973 (.CO(inst_cellmath__63__W0[7]), .S(inst_cellmath__63__W1[6]), .A(N6117), .B(N6529), .CI(N6495));
ADDHX1 inst_cellmath__63_0_I1974 (.CO(N6574), .S(N6388), .A(N6186), .B(N6328));
ADDFX1 inst_cellmath__63_0_I1975 (.CO(N6085), .S(N5898), .A(N6213), .B(N6268), .CI(N6128));
ADDFX1 inst_cellmath__63_0_I1976 (.CO(N6464), .S(N6273), .A(N6154), .B(N6240), .CI(N6295));
ADDFX1 inst_cellmath__63_0_I1977 (.CO(N5979), .S(N5791), .A(N5931), .B(N6417), .CI(N6388));
ADDFX1 inst_cellmath__63_0_I1978 (.CO(N6357), .S(N6164), .A(N6306), .B(N5898), .CI(N6273));
ADDFX1 inst_cellmath__63_0_I1979 (.CO(inst_cellmath__63__W0[8]), .S(inst_cellmath__63__W1[7]), .A(N5791), .B(N5821), .CI(N6164));
ADDHX1 inst_cellmath__63_0_I1980 (.CO(N6244), .S(N6055), .A(N5730), .B(N5867));
ADDFX1 inst_cellmath__63_0_I1981 (.CO(N5758), .S(N6433), .A(N5754), .B(N5813), .CI(N6503));
ADDFX1 inst_cellmath__63_0_I1982 (.CO(N6136), .S(N5948), .A(N6535), .B(N5785), .CI(N6560));
ADDFX1 inst_cellmath__63_0_I1983 (.CO(N6513), .S(N6324), .A(N6574), .B(N5841), .CI(N6055));
ADDFX1 inst_cellmath__63_0_I1984 (.CO(N6026), .S(N5839), .A(N6464), .B(N6085), .CI(N6433));
ADDFX1 inst_cellmath__63_0_I1985 (.CO(N6404), .S(N6212), .A(N5979), .B(N5948), .CI(N6324));
ADDFX1 inst_cellmath__63_0_I1986 (.CO(inst_cellmath__63__W0[9]), .S(inst_cellmath__63__W1[8]), .A(N5839), .B(N6357), .CI(N6212));
ADDHX1 inst_cellmath__63_0_I1987 (.CO(N6289), .S(N6101), .A(N6132), .B(N6270));
ADDFX1 inst_cellmath__63_0_I1988 (.CO(N5806), .S(N6480), .A(N6018), .B(N6216), .CI(N6042));
ADDFX1 inst_cellmath__63_0_I1989 (.CO(N6181), .S(N5993), .A(N6157), .B(N6189), .CI(N6073));
ADDFX1 inst_cellmath__63_0_I1990 (.CO(N6557), .S(N6370), .A(N6243), .B(N6100), .CI(N6244));
ADDFX1 inst_cellmath__63_0_I1991 (.CO(N6069), .S(N5880), .A(N5758), .B(N6101), .CI(N6136));
ADDFX1 inst_cellmath__63_0_I1992 (.CO(N6447), .S(N6255), .A(N6480), .B(N5993), .CI(N6513));
ADDFX1 inst_cellmath__63_0_I1993 (.CO(N5960), .S(N5772), .A(N6026), .B(N6370), .CI(N5880));
ADDFX1 inst_cellmath__63_0_I1994 (.CO(inst_cellmath__63__W0[10]), .S(inst_cellmath__63__W1[9]), .A(N6255), .B(N6404), .CI(N5772));
ADDHX1 inst_cellmath__63_0_I1995 (.CO(N5849), .S(N6524), .A(N6538), .B(N5815));
ADDFX1 inst_cellmath__63_0_I1996 (.CO(N6224), .S(N6036), .A(N6422), .B(N5756), .CI(N6452));
ADDFX1 inst_cellmath__63_0_I1997 (.CO(N5739), .S(N6413), .A(N6562), .B(N6398), .CI(N6481));
ADDFX1 inst_cellmath__63_0_I1998 (.CO(N6115), .S(N5928), .A(N6509), .B(N5733), .CI(N5787));
ADDFX1 inst_cellmath__63_0_I1999 (.CO(N6492), .S(N6302), .A(N6524), .B(N6289), .CI(N5806));
ADDFX1 inst_cellmath__63_0_I2000 (.CO(N6007), .S(N5818), .A(N6413), .B(N6181), .CI(N6036));
ADDFX1 inst_cellmath__63_0_I2001 (.CO(N6386), .S(N6195), .A(N5928), .B(N6557), .CI(N6069));
ADDFX1 inst_cellmath__63_0_I2002 (.CO(N5895), .S(N6571), .A(N6447), .B(N6302), .CI(N5818));
ADDFX1 inst_cellmath__63_0_I2003 (.CO(inst_cellmath__63__W0[11]), .S(inst_cellmath__63__W1[10]), .A(N5960), .B(N6195), .CI(N6571));
ADDHX1 inst_cellmath__63_0_I2004 (.CO(N5789), .S(N6462), .A(N6076), .B(N6219));
ADDFX1 inst_cellmath__63_0_I2005 (.CO(N6161), .S(N5976), .A(N5964), .B(N6158), .CI(N5994));
ADDFX1 inst_cellmath__63_0_I2006 (.CO(N6542), .S(N6352), .A(N6103), .B(N5935), .CI(N6022));
ADDFX1 inst_cellmath__63_0_I2007 (.CO(N6051), .S(N5864), .A(N6047), .B(N6134), .CI(N6191));
ADDFX1 inst_cellmath__63_0_I2008 (.CO(N6428), .S(N6239), .A(N5849), .B(N5906), .CI(N6462));
ADDFX1 inst_cellmath__63_0_I2009 (.CO(N5943), .S(N5753), .A(N6224), .B(N5739), .CI(N6115));
ADDFX1 inst_cellmath__63_0_I2010 (.CO(N6320), .S(N6131), .A(N5976), .B(N6352), .CI(N5864));
ADDFX1 inst_cellmath__63_0_I2011 (.CO(N5834), .S(N6508), .A(N6239), .B(N6492), .CI(N6007));
ADDFX1 inst_cellmath__63_0_I2012 (.CO(N6208), .S(N6021), .A(N6386), .B(N5753), .CI(N6131));
ADDFX1 inst_cellmath__63_0_I2013 (.CO(inst_cellmath__63__W0[12]), .S(inst_cellmath__63__W1[11]), .A(N5895), .B(N6508), .CI(N6021));
ADDHX1 inst_cellmath__63_0_I2014 (.CO(N6096), .S(N5911), .A(N6484), .B(N5759));
ADDFX1 inst_cellmath__63_0_I2015 (.CO(N6476), .S(N6284), .A(N6369), .B(N6564), .CI(N6400));
ADDFX1 inst_cellmath__63_0_I2016 (.CO(N5988), .S(N5801), .A(N6512), .B(N6341), .CI(N6424));
ADDFX1 inst_cellmath__63_0_I2017 (.CO(N6365), .S(N6176), .A(N6455), .B(N6540), .CI(N6311));
ADDFX1 inst_cellmath__63_0_I2018 (.CO(N5876), .S(N6552), .A(N5735), .B(N6282), .CI(N5789));
ADDFX1 inst_cellmath__63_0_I2019 (.CO(N6251), .S(N6064), .A(N6542), .B(N5911), .CI(N6161));
ADDFX1 inst_cellmath__63_0_I2020 (.CO(N5767), .S(N6441), .A(N5801), .B(N6051), .CI(N6284));
ADDFX1 inst_cellmath__63_0_I2021 (.CO(N6142), .S(N5955), .A(N6428), .B(N6176), .CI(N5943));
ADDFX1 inst_cellmath__63_0_I2022 (.CO(N6521), .S(N6332), .A(N6064), .B(N6552), .CI(N6320));
ADDFX1 inst_cellmath__63_0_I2023 (.CO(N6032), .S(N5846), .A(N5834), .B(N6441), .CI(N5955));
ADDFX1 inst_cellmath__63_0_I2024 (.CO(inst_cellmath__63__W0[13]), .S(inst_cellmath__63__W1[12]), .A(N6332), .B(N6208), .CI(N5846));
ADDHX1 inst_cellmath__63_0_I2025 (.CO(N5924), .S(N5737), .A(N6024), .B(N6162));
ADDFX1 inst_cellmath__63_0_I2026 (.CO(N6298), .S(N6111), .A(N5799), .B(N6106), .CI(N5939));
ADDFX1 inst_cellmath__63_0_I2027 (.CO(N5816), .S(N6490), .A(N5912), .B(N5881), .CI(N5966));
ADDFX1 inst_cellmath__63_0_I2028 (.CO(N6192), .S(N6004), .A(N6049), .B(N6079), .CI(N5997));
ADDFX1 inst_cellmath__63_0_I2029 (.CO(N6566), .S(N6382), .A(N6138), .B(N5826), .CI(N5853));
ADDFX1 inst_cellmath__63_0_I2030 (.CO(N6080), .S(N5891), .A(N5737), .B(N6096), .CI(N6476));
ADDFX1 inst_cellmath__63_0_I2031 (.CO(N6458), .S(N6267), .A(N6365), .B(N5988), .CI(N6490));
ADDFX1 inst_cellmath__63_0_I2032 (.CO(N5970), .S(N5784), .A(N6004), .B(N6111), .CI(N5876));
ADDFX1 inst_cellmath__63_0_I2033 (.CO(N6347), .S(N6156), .A(N6251), .B(N6382), .CI(N5767));
ADDFX1 inst_cellmath__63_0_I2034 (.CO(N5859), .S(N6537), .A(N6267), .B(N5891), .CI(N6142));
ADDFX1 inst_cellmath__63_0_I2035 (.CO(N6233), .S(N6046), .A(N6521), .B(N5784), .CI(N6156));
ADDFX1 inst_cellmath__63_0_I2036 (.CO(inst_cellmath__63__W0[14]), .S(inst_cellmath__63__W1[13]), .A(N6032), .B(N6537), .CI(N6046));
ADDHX1 inst_cellmath__63_0_I2037 (.CO(N6126), .S(N5938), .A(N6172), .B(N6201));
ADDFX1 inst_cellmath__63_0_I2038 (.CO(N6502), .S(N6315), .A(N6515), .B(N6425), .CI(N6344));
ADDFX1 inst_cellmath__63_0_I2039 (.CO(N6016), .S(N5829), .A(N6316), .B(N6285), .CI(N6373));
ADDFX1 inst_cellmath__63_0_I2040 (.CO(N6396), .S(N6204), .A(N6457), .B(N6486), .CI(N6401));
ADDFX1 inst_cellmath__63_0_I2041 (.CO(N5905), .S(N5723), .A(N6567), .B(N6227), .CI(N6256));
ADDFX1 inst_cellmath__63_0_I2042 (.CO(N6280), .S(N6091), .A(N5924), .B(N6543), .CI(N5938));
ADDFX1 inst_cellmath__63_0_I2043 (.CO(N5797), .S(N6472), .A(N6192), .B(N5816), .CI(N6298));
ADDFX1 inst_cellmath__63_0_I2044 (.CO(N6171), .S(N5984), .A(N5829), .B(N6566), .CI(N6204));
ADDFX1 inst_cellmath__63_0_I2045 (.CO(N6548), .S(N6362), .A(N5723), .B(N6315), .CI(N6080));
ADDFX1 inst_cellmath__63_0_I2046 (.CO(N6060), .S(N5872), .A(N6458), .B(N6091), .CI(N6472));
ADDFX1 inst_cellmath__63_0_I2047 (.CO(N6437), .S(N6248), .A(N5984), .B(N5970), .CI(N6362));
ADDFX1 inst_cellmath__63_0_I2048 (.CO(N5952), .S(N5764), .A(N5872), .B(N6347), .CI(N5859));
ADDFX1 inst_cellmath__63_0_I2049 (.CO(inst_cellmath__63__W0[15]), .S(inst_cellmath__63__W1[14]), .A(N6248), .B(N6233), .CI(N5764));
XNOR2X1 inst_cellmath__63_0_I2050 (.Y(N6518), .A(N6108), .B(N6550));
OR2XL inst_cellmath__63_0_I2051 (.Y(N5843), .A(N6108), .B(N6550));
ADDFX1 inst_cellmath__63_0_I2052 (.CO(N5736), .S(N6410), .A(N5968), .B(N6580), .CI(N5883));
ADDFX1 inst_cellmath__63_0_I2053 (.CO(N6107), .S(N5920), .A(N5743), .B(N6052), .CI(N5915));
ADDFX1 inst_cellmath__63_0_I2054 (.CO(N6487), .S(N6296), .A(N5856), .B(N5830), .CI(N6000));
ADDFX1 inst_cellmath__63_0_I2055 (.CO(N6001), .S(N5812), .A(N5941), .B(N6027), .CI(N5802));
ADDFX1 inst_cellmath__63_0_I2056 (.CO(N6377), .S(N6188), .A(N6081), .B(N5771), .CI(N6126));
ADDFX1 inst_cellmath__63_0_I2057 (.CO(N5887), .S(N6563), .A(N6016), .B(N6518), .CI(N6396));
ADDFX1 inst_cellmath__63_0_I2058 (.CO(N6263), .S(N6075), .A(N5905), .B(N6502), .CI(N6296));
ADDFX1 inst_cellmath__63_0_I2059 (.CO(N5779), .S(N6454), .A(N6410), .B(N5920), .CI(N5812));
ADDFX1 inst_cellmath__63_0_I2060 (.CO(N6152), .S(N5967), .A(N6188), .B(N6280), .CI(N5797));
ADDFX1 inst_cellmath__63_0_I2061 (.CO(N6532), .S(N6343), .A(N6171), .B(N6563), .CI(N6075));
ADDFX1 inst_cellmath__63_0_I2062 (.CO(N6040), .S(N5855), .A(N6454), .B(N6548), .CI(N6060));
ADDFX1 inst_cellmath__63_0_I2063 (.CO(N6420), .S(N6230), .A(N6343), .B(N5967), .CI(N6437));
ADDFX1 inst_cellmath__63_0_I2064 (.CO(inst_cellmath__63__W0[16]), .S(inst_cellmath__63__W1[15]), .A(N5952), .B(N5855), .CI(N6230));
ADDFX1 inst_cellmath__63_0_I2065 (.CO(N6309), .S(N6120), .A(N6488), .B(N6062), .CI(N6088));
ADDFX1 inst_cellmath__63_0_I2066 (.CO(N5824), .S(N6498), .A(N6376), .B(N6118), .CI(N6287));
ADDFX1 inst_cellmath__63_0_I2067 (.CO(N6199), .S(N6011), .A(N6146), .B(N6459), .CI(N6318));
ADDFX1 inst_cellmath__63_0_I2068 (.CO(N6577), .S(N6391), .A(N6259), .B(N6229), .CI(N6406));
ADDFX1 inst_cellmath__63_0_I2069 (.CO(N6086), .S(N5901), .A(N6346), .B(N6429), .CI(N6205));
ADDFX1 inst_cellmath__63_0_I2070 (.CO(N6467), .S(N6275), .A(N5843), .B(N6177), .CI(N6487));
ADDFX1 inst_cellmath__63_0_I2071 (.CO(N5981), .S(N5793), .A(N5736), .B(N6107), .CI(N6120));
ADDFX1 inst_cellmath__63_0_I2072 (.CO(N6359), .S(N6167), .A(N6377), .B(N6001), .CI(N6498));
ADDFX1 inst_cellmath__63_0_I2073 (.CO(N5870), .S(N6547), .A(N6011), .B(N6391), .CI(N5901));
ADDFX1 inst_cellmath__63_0_I2074 (.CO(N6246), .S(N6057), .A(N6263), .B(N5887), .CI(N6275));
ADDFX1 inst_cellmath__63_0_I2075 (.CO(N5760), .S(N6435), .A(N5779), .B(N5793), .CI(N6167));
ADDFX1 inst_cellmath__63_0_I2076 (.CO(N6139), .S(N5950), .A(N6547), .B(N6152), .CI(N6532));
ADDFX1 inst_cellmath__63_0_I2077 (.CO(N6516), .S(N6327), .A(N6040), .B(N6057), .CI(N6435));
ADDFX1 inst_cellmath__63_0_I2078 (.CO(inst_cellmath__63__W0[17]), .S(inst_cellmath__63__W1[16]), .A(N6420), .B(N5950), .CI(N6327));
ADDFX1 inst_cellmath__63_0_I2079 (.CO(N6407), .S(N6215), .A(N6002), .B(N6438), .CI(N6469));
ADDFX1 inst_cellmath__63_0_I2080 (.CO(N5917), .S(N5732), .A(N6525), .B(N6494), .CI(N5916));
ADDFX1 inst_cellmath__63_0_I2081 (.CO(N6292), .S(N6102), .A(N6553), .B(N5775), .CI(N5831));
ADDFX1 inst_cellmath__63_0_I2082 (.CO(N5809), .S(N6483), .A(N5804), .B(N5972), .CI(N5858));
ADDFX1 inst_cellmath__63_0_I2083 (.CO(N6184), .S(N5996), .A(N5886), .B(N5944), .CI(N5745));
ADDFX1 inst_cellmath__63_0_I2084 (.CO(N6559), .S(N6372), .A(N6215), .B(N5724), .CI(N6309));
ADDFX1 inst_cellmath__63_0_I2085 (.CO(N6072), .S(N5882), .A(N6199), .B(N6577), .CI(N5824));
ADDFX1 inst_cellmath__63_0_I2086 (.CO(N6450), .S(N6258), .A(N5732), .B(N6086), .CI(N6483));
ADDFX1 inst_cellmath__63_0_I2087 (.CO(N5962), .S(N5774), .A(N5996), .B(N6102), .CI(N6467));
ADDFX1 inst_cellmath__63_0_I2088 (.CO(N6339), .S(N6147), .A(N6372), .B(N5981), .CI(N6359));
ADDFX1 inst_cellmath__63_0_I2089 (.CO(N5851), .S(N6527), .A(N5870), .B(N5882), .CI(N6258));
ADDFX1 inst_cellmath__63_0_I2090 (.CO(N6226), .S(N6037), .A(N6246), .B(N5774), .CI(N6147));
ADDFX1 inst_cellmath__63_0_I2091 (.CO(N5741), .S(N6415), .A(N6527), .B(N5760), .CI(N6139));
ADDFX1 inst_cellmath__63_0_I2092 (.CO(inst_cellmath__63__W0[18]), .S(inst_cellmath__63__W1[17]), .A(N6516), .B(N6037), .CI(N6415));
INVXL inst_cellmath__63_0_I2093 (.Y(N5922), .A(N6301));
ADDFX1 inst_cellmath__63_0_I2094 (.CO(N6493), .S(N6303), .A(N6378), .B(N5982), .CI(N5922));
ADDFX1 inst_cellmath__63_0_I2095 (.CO(N6387), .S(N6196), .A(N6034), .B(N6009), .CI(N6065));
ADDFX1 inst_cellmath__63_0_I2096 (.CO(N5896), .S(N6572), .A(N6180), .B(N6321), .CI(N6232));
ADDFX1 inst_cellmath__63_0_I2097 (.CO(N6272), .S(N6084), .A(N6092), .B(N6348), .CI(N6121));
ADDFX1 inst_cellmath__63_0_I2098 (.CO(N5790), .S(N6463), .A(N6262), .B(N6206), .CI(N6290));
ADDFX1 inst_cellmath__63_0_I2099 (.CO(N6163), .S(N5978), .A(N6148), .B(N6407), .CI(N6303));
ADDFX1 inst_cellmath__63_0_I2100 (.CO(N6545), .S(N6354), .A(N5809), .B(N5917), .CI(N6292));
ADDFX1 inst_cellmath__63_0_I2101 (.CO(N6053), .S(N5866), .A(N6184), .B(N6196), .CI(N6572));
ADDFX1 inst_cellmath__63_0_I2102 (.CO(N6430), .S(N6242), .A(N6084), .B(N6463), .CI(N6559));
ADDFX1 inst_cellmath__63_0_I2103 (.CO(N5946), .S(N5755), .A(N5978), .B(N6072), .CI(N6450));
ADDFX1 inst_cellmath__63_0_I2104 (.CO(N6322), .S(N6133), .A(N5962), .B(N6354), .CI(N5866));
ADDFX1 inst_cellmath__63_0_I2105 (.CO(N5836), .S(N6511), .A(N6339), .B(N6242), .CI(N5755));
ADDFX1 inst_cellmath__63_0_I2106 (.CO(N6211), .S(N6023), .A(N6133), .B(N5851), .CI(N6226));
ADDFX1 inst_cellmath__63_0_I2107 (.CO(inst_cellmath__63__W0[19]), .S(inst_cellmath__63__W1[18]), .A(N5741), .B(N6511), .CI(N6023));
ADDFX1 inst_cellmath__63_0_I2108 (.CO(N6098), .S(N5914), .A(N6301), .B(N6570), .CI(N6389));
ADDFX1 inst_cellmath__63_0_I2109 (.CO(N6479), .S(N6286), .A(N6414), .B(N5888), .CI(N5914));
ADDFX1 inst_cellmath__63_0_I2110 (.CO(N5990), .S(N5803), .A(N6473), .B(N6442), .CI(N5860));
ADDFX1 inst_cellmath__63_0_I2111 (.CO(N6367), .S(N6179), .A(N6493), .B(N5726), .CI(N5778));
ADDFX1 inst_cellmath__63_0_I2112 (.CO(N5879), .S(N6554), .A(N6497), .B(N5747), .CI(N6528));
ADDFX1 inst_cellmath__63_0_I2113 (.CO(N6253), .S(N6066), .A(N5835), .B(N5808), .CI(N6555));
ADDFX1 inst_cellmath__63_0_I2114 (.CO(N5769), .S(N6444), .A(N6286), .B(N6387), .CI(N5896));
ADDFX1 inst_cellmath__63_0_I2115 (.CO(N6145), .S(N5957), .A(N6272), .B(N5790), .CI(N5803));
ADDFX1 inst_cellmath__63_0_I2116 (.CO(N6523), .S(N6334), .A(N6163), .B(N6554), .CI(N6066));
ADDFX1 inst_cellmath__63_0_I2117 (.CO(N6033), .S(N5847), .A(N6545), .B(N6179), .CI(N6053));
ADDFX1 inst_cellmath__63_0_I2118 (.CO(N6412), .S(N6222), .A(N6430), .B(N6444), .CI(N5957));
ADDFX1 inst_cellmath__63_0_I2119 (.CO(N5927), .S(N5738), .A(N5946), .B(N6334), .CI(N5847));
ADDFX1 inst_cellmath__63_0_I2120 (.CO(N6299), .S(N6112), .A(N6222), .B(N6322), .CI(N5836));
ADDFX1 inst_cellmath__63_0_I2121 (.CO(inst_cellmath__63__W0[20]), .S(inst_cellmath__63__W1[19]), .A(N6211), .B(N5738), .CI(N6112));
ADDFX1 inst_cellmath__63_0_I2122 (.CO(N6194), .S(N6005), .A(N5929), .B(N5975), .CI(N6098));
ADDFX1 inst_cellmath__63_0_I2123 (.CO(N6568), .S(N6384), .A(N5956), .B(N6264), .CI(N5985));
ADDFX1 inst_cellmath__63_0_I2124 (.CO(N6082), .S(N5894), .A(N6124), .B(N6012), .CI(N6183));
ADDFX1 inst_cellmath__63_0_I2125 (.CO(N6461), .S(N6269), .A(N6038), .B(N6151), .CI(N6067));
ADDFX1 inst_cellmath__63_0_I2126 (.CO(N5973), .S(N5786), .A(N6235), .B(N6209), .CI(N6093));
ADDFX1 inst_cellmath__63_0_I2127 (.CO(N6350), .S(N6160), .A(N6005), .B(N6479), .CI(N5990));
ADDFX1 inst_cellmath__63_0_I2128 (.CO(N5863), .S(N6539), .A(N6384), .B(N5879), .CI(N6253));
ADDFX1 inst_cellmath__63_0_I2129 (.CO(N6236), .S(N6048), .A(N5894), .B(N6367), .CI(N6269));
ADDFX1 inst_cellmath__63_0_I2130 (.CO(N5751), .S(N6427), .A(N5769), .B(N5786), .CI(N6145));
ADDFX1 inst_cellmath__63_0_I2131 (.CO(N6130), .S(N5940), .A(N6523), .B(N6160), .CI(N6539));
ADDFX1 inst_cellmath__63_0_I2132 (.CO(N6505), .S(N6317), .A(N6033), .B(N6048), .CI(N6427));
ADDFX1 inst_cellmath__63_0_I2133 (.CO(N6019), .S(N5833), .A(N5940), .B(N6412), .CI(N5927));
ADDFX1 inst_cellmath__63_0_I2134 (.CO(inst_cellmath__63__W0[21]), .S(inst_cellmath__63__W1[20]), .A(N6299), .B(N6317), .CI(N5833));
ADDFX1 inst_cellmath__63_0_I2135 (.CO(N5908), .S(N5725), .A(N6333), .B(N2876), .CI(N5780));
ADDFX1 inst_cellmath__63_0_I2136 (.CO(N6283), .S(N6095), .A(N6392), .B(N6361), .CI(N6416));
ADDFX1 inst_cellmath__63_0_I2137 (.CO(N5800), .S(N6474), .A(N6531), .B(N6194), .CI(N5728));
ADDFX1 inst_cellmath__63_0_I2138 (.CO(N6174), .S(N5986), .A(N6445), .B(N6558), .CI(N6475));
ADDFX1 inst_cellmath__63_0_I2139 (.CO(N6551), .S(N6364), .A(N6501), .B(N5749), .CI(N5725));
ADDFX1 inst_cellmath__63_0_I2140 (.CO(N6063), .S(N5874), .A(N6082), .B(N6568), .CI(N6461));
ADDFX1 inst_cellmath__63_0_I2141 (.CO(N6439), .S(N6249), .A(N5973), .B(N6095), .CI(N6474));
ADDFX1 inst_cellmath__63_0_I2142 (.CO(N5954), .S(N5766), .A(N6350), .B(N5986), .CI(N6364));
ADDFX1 inst_cellmath__63_0_I2143 (.CO(N6331), .S(N6141), .A(N5874), .B(N5863), .CI(N6236));
ADDFX1 inst_cellmath__63_0_I2144 (.CO(N5844), .S(N6519), .A(N5751), .B(N6249), .CI(N5766));
ADDFX1 inst_cellmath__63_0_I2145 (.CO(N6220), .S(N6031), .A(N6141), .B(N6130), .CI(N6505));
ADDFX1 inst_cellmath__63_0_I2146 (.CO(inst_cellmath__63__W0[22]), .S(inst_cellmath__63__W1[21]), .A(N6019), .B(N6519), .CI(N6031));
ADDFX1 inst_cellmath__63_0_I2147 (.CO(N6109), .S(N5923), .A(N5873), .B(N11660), .CI(N6153));
ADDFX1 inst_cellmath__63_0_I2148 (.CO(N6489), .S(N6297), .A(N5930), .B(N5900), .CI(N5958));
ADDFX1 inst_cellmath__63_0_I2149 (.CO(N6003), .S(N5814), .A(N5908), .B(N6071), .CI(N6127));
ADDFX1 inst_cellmath__63_0_I2150 (.CO(N6380), .S(N6190), .A(N5987), .B(N6097), .CI(N6014));
ADDFX1 inst_cellmath__63_0_I2151 (.CO(N5890), .S(N6565), .A(N5923), .B(N6039), .CI(N6283));
ADDFX1 inst_cellmath__63_0_I2152 (.CO(N6266), .S(N6078), .A(N6174), .B(N5800), .CI(N6297));
ADDFX1 inst_cellmath__63_0_I2153 (.CO(N5782), .S(N6456), .A(N6190), .B(N6551), .CI(N5814));
ADDFX1 inst_cellmath__63_0_I2154 (.CO(N6155), .S(N5969), .A(N6565), .B(N6063), .CI(N6439));
ADDFX1 inst_cellmath__63_0_I2155 (.CO(N6536), .S(N6345), .A(N5954), .B(N6078), .CI(N6456));
ADDFX1 inst_cellmath__63_0_I2156 (.CO(N6043), .S(N5857), .A(N5969), .B(N6331), .CI(N5844));
ADDFX1 inst_cellmath__63_0_I2157 (.CO(inst_cellmath__63__W0[23]), .S(inst_cellmath__63__W1[22]), .A(N6220), .B(N6345), .CI(N5857));
ADDFX1 inst_cellmath__63_0_I2158 (.CO(N5937), .S(N5746), .A(N6276), .B(N11669), .CI(N6534));
ADDFX1 inst_cellmath__63_0_I2159 (.CO(N6312), .S(N6123), .A(N6335), .B(N6304), .CI(N6363));
ADDFX1 inst_cellmath__63_0_I2160 (.CO(N5827), .S(N6500), .A(N6477), .B(N6109), .CI(N6394));
ADDFX1 inst_cellmath__63_0_I2161 (.CO(N6203), .S(N6013), .A(N6419), .B(N6504), .CI(N6449));
ADDFX1 inst_cellmath__63_0_I2162 (.CO(N6581), .S(N6393), .A(N6489), .B(N5746), .CI(N6380));
ADDFX1 inst_cellmath__63_0_I2163 (.CO(N6089), .S(N5903), .A(N6123), .B(N6003), .CI(N6500));
ADDFX1 inst_cellmath__63_0_I2164 (.CO(N6471), .S(N6277), .A(N6013), .B(N5890), .CI(N6266));
ADDFX1 inst_cellmath__63_0_I2165 (.CO(N5983), .S(N5794), .A(N5782), .B(N6393), .CI(N5903));
ADDFX1 inst_cellmath__63_0_I2166 (.CO(N6360), .S(N6169), .A(N6277), .B(N6155), .CI(N6536));
ADDFX1 inst_cellmath__63_0_I2167 (.CO(inst_cellmath__63__W0[24]), .S(inst_cellmath__63__W1[23]), .A(N6043), .B(N5794), .CI(N6169));
ADDFX1 inst_cellmath__63_0_I2168 (.CO(N6247), .S(N6058), .A(N5820), .B(N2773), .CI(N6041));
ADDFX1 inst_cellmath__63_0_I2169 (.CO(N5762), .S(N6436), .A(N5875), .B(N5848), .CI(N5904));
ADDFX1 inst_cellmath__63_0_I2170 (.CO(N6140), .S(N5951), .A(N6017), .B(N5937), .CI(N5933));
ADDFX1 inst_cellmath__63_0_I2171 (.CO(N6517), .S(N6329), .A(N5989), .B(N5961), .CI(N6058));
ADDFX1 inst_cellmath__63_0_I2172 (.CO(N6030), .S(N5842), .A(N5827), .B(N6312), .CI(N6436));
ADDFX1 inst_cellmath__63_0_I2173 (.CO(N6409), .S(N6218), .A(N5951), .B(N6203), .CI(N6329));
ADDFX1 inst_cellmath__63_0_I2174 (.CO(N5919), .S(N5734), .A(N6089), .B(N6581), .CI(N5842));
ADDFX1 inst_cellmath__63_0_I2175 (.CO(N6294), .S(N6105), .A(N6218), .B(N6471), .CI(N5983));
ADDFX1 inst_cellmath__63_0_I2176 (.CO(inst_cellmath__63__W0[25]), .S(inst_cellmath__63__W1[24]), .A(N6360), .B(N5734), .CI(N6105));
ADDFX1 inst_cellmath__63_0_I2177 (.CO(N6187), .S(N5999), .A(N6223), .B(N11688), .CI(N6421));
ADDFX1 inst_cellmath__63_0_I2178 (.CO(N6561), .S(N6375), .A(N6278), .B(N6250), .CI(N6308));
ADDFX1 inst_cellmath__63_0_I2179 (.CO(N6074), .S(N5885), .A(N6338), .B(N6247), .CI(N6366));
ADDFX1 inst_cellmath__63_0_I2180 (.CO(N6453), .S(N6261), .A(N5999), .B(N6397), .CI(N5762));
ADDFX1 inst_cellmath__63_0_I2181 (.CO(N5965), .S(N5777), .A(N6375), .B(N6140), .CI(N6517));
ADDFX1 inst_cellmath__63_0_I2182 (.CO(N6342), .S(N6150), .A(N6261), .B(N5885), .CI(N6030));
ADDFX1 inst_cellmath__63_0_I2183 (.CO(N5854), .S(N6530), .A(N6409), .B(N5777), .CI(N5919));
ADDFX1 inst_cellmath__63_0_I2184 (.CO(inst_cellmath__63__W0[26]), .S(inst_cellmath__63__W1[25]), .A(N6294), .B(N6150), .CI(N6530));
ADDFX1 inst_cellmath__63_0_I2185 (.CO(N5744), .S(N6418), .A(N5765), .B(N11697), .CI(N5795));
ADDFX1 inst_cellmath__63_0_I2186 (.CO(N6119), .S(N5932), .A(N5823), .B(N5934), .CI(N5850));
ADDFX1 inst_cellmath__63_0_I2187 (.CO(N6496), .S(N6307), .A(N5877), .B(N6187), .CI(N5907));
ADDFX1 inst_cellmath__63_0_I2188 (.CO(N6010), .S(N5822), .A(N6561), .B(N6418), .CI(N6074));
ADDFX1 inst_cellmath__63_0_I2189 (.CO(N6390), .S(N6197), .A(N6307), .B(N5932), .CI(N6453));
ADDFX1 inst_cellmath__63_0_I2190 (.CO(N5899), .S(N6575), .A(N5822), .B(N5965), .CI(N6197));
ADDFX1 inst_cellmath__63_0_I2191 (.CO(inst_cellmath__63__W1[27]), .S(inst_cellmath__63__W1[26]), .A(N5854), .B(N6342), .CI(N6575));
ADDFX1 inst_cellmath__63_0_I2192 (.CO(N5792), .S(N6465), .A(N6170), .B(N11706), .CI(N6310));
ADDFX1 inst_cellmath__63_0_I2193 (.CO(N6165), .S(N5980), .A(N6225), .B(N6198), .CI(N6252));
ADDFX1 inst_cellmath__63_0_I2194 (.CO(N6546), .S(N6358), .A(N5744), .B(N6281), .CI(N6465));
ADDFX1 inst_cellmath__63_0_I2195 (.CO(N6056), .S(N5869), .A(N6496), .B(N6119), .CI(N5980));
ADDFX1 inst_cellmath__63_0_I2196 (.CO(N6434), .S(N6245), .A(N6010), .B(N6358), .CI(N5869));
ADDFX1 inst_cellmath__63_0_I2197 (.CO(inst_cellmath__63__W1[28]), .S(inst_cellmath__63__W0[27]), .A(N6245), .B(N6390), .CI(N5899));
ADDFX1 inst_cellmath__63_0_I2198 (.CO(N6326), .S(N6137), .A(N6576), .B(N11708), .CI(N5825));
ADDFX1 inst_cellmath__63_0_I2199 (.CO(N5840), .S(N6514), .A(N5768), .B(N5740), .CI(N5798));
ADDFX1 inst_cellmath__63_0_I2200 (.CO(N6214), .S(N6028), .A(N6137), .B(N5792), .CI(N6165));
ADDFX1 inst_cellmath__63_0_I2201 (.CO(N5731), .S(N6405), .A(N6546), .B(N6514), .CI(N6028));
ADDFX1 inst_cellmath__63_0_I2202 (.CO(inst_cellmath__63__W1[29]), .S(inst_cellmath__63__W0[28]), .A(N6405), .B(N6056), .CI(N6434));
ADDFX1 inst_cellmath__63_0_I2203 (.CO(N6482), .S(N6291), .A(N6116), .B(N11719), .CI(N6200));
ADDFX1 inst_cellmath__63_0_I2204 (.CO(N5995), .S(N5807), .A(N6173), .B(N6143), .CI(N6326));
ADDFX1 inst_cellmath__63_0_I2205 (.CO(N6371), .S(N6182), .A(N5840), .B(N6291), .CI(N5807));
ADDFX1 inst_cellmath__63_0_I2206 (.CO(inst_cellmath__63__W1[30]), .S(inst_cellmath__63__W0[29]), .A(N6182), .B(N6214), .CI(N5731));
ADDFX1 inst_cellmath__63_0_I2207 (.CO(N6257), .S(N6070), .A(N6522), .B(N11728), .CI(N6579));
ADDFX1 inst_cellmath__63_0_I2208 (.CO(N5773), .S(N6448), .A(N6482), .B(N6549), .CI(N6070));
ADDFX1 inst_cellmath__63_0_I2209 (.CO(inst_cellmath__63__W1[31]), .S(inst_cellmath__63__W0[30]), .A(N6448), .B(N5995), .CI(N6371));
ADDFX1 inst_cellmath__63_0_I2210 (.CO(N6526), .S(N6337), .A(N6061), .B(N2705), .CI(N6087));
ADDFX1 inst_cellmath__63_0_I2211 (.CO(inst_cellmath__63__W1[32]), .S(inst_cellmath__63__W0[31]), .A(N6337), .B(N6257), .CI(N5773));
ADDFX1 inst_cellmath__63_0_I2212 (.CO(inst_cellmath__63__W1[33]), .S(inst_cellmath__63__W0[32]), .A(N6468), .B(N2777), .CI(N6526));
ADDHX1 cynw_cm_float_rcp_I2213 (.CO(N7618), .S(N7487), .A(N477), .B(inst_cellmath__63__W0[15]));
XNOR2X1 cynw_cm_float_rcp_I2214 (.Y(N7757), .A(N478), .B(inst_cellmath__63__W0[16]));
OR2XL cynw_cm_float_rcp_I2215 (.Y(N7890), .A(N478), .B(inst_cellmath__63__W0[16]));
ADDHX1 cynw_cm_float_rcp_I2216 (.CO(N7806), .S(N7675), .A(inst_cellmath__63__W1[16]), .B(inst_cellmath__62__W0[16]));
ADDFX1 cynw_cm_float_rcp_I2217 (.CO(N7457), .S(N7945), .A(inst_cellmath__63__W0[17]), .B(N479), .CI(inst_cellmath__63__W1[17]));
ADDHX1 cynw_cm_float_rcp_I2218 (.CO(N7730), .S(N7597), .A(inst_cellmath__62__W0[17]), .B(inst_cellmath__62__W1[17]));
ADDFX1 cynw_cm_float_rcp_I2219 (.CO(N8001), .S(N7864), .A(inst_cellmath__63__W0[18]), .B(N480), .CI(inst_cellmath__63__W1[18]));
ADDHX1 cynw_cm_float_rcp_I2220 (.CO(N7649), .S(N7520), .A(inst_cellmath__62__W0[18]), .B(inst_cellmath__62__W1[18]));
ADDFX1 cynw_cm_float_rcp_I2221 (.CO(N7924), .S(N7787), .A(inst_cellmath__63__W0[19]), .B(N481), .CI(inst_cellmath__63__W1[19]));
ADDHX1 cynw_cm_float_rcp_I2222 (.CO(N7575), .S(N7434), .A(inst_cellmath__62__W0[19]), .B(inst_cellmath__62__W1[19]));
ADDFX1 cynw_cm_float_rcp_I2223 (.CO(N7838), .S(N7709), .A(inst_cellmath__63__W0[20]), .B(N482), .CI(inst_cellmath__63__W1[20]));
ADDHX1 cynw_cm_float_rcp_I2224 (.CO(N7497), .S(N7980), .A(inst_cellmath__62__W0[20]), .B(inst_cellmath__62__W1[20]));
ADDFX1 cynw_cm_float_rcp_I2225 (.CO(N7767), .S(N7627), .A(inst_cellmath__63__W0[21]), .B(N483), .CI(inst_cellmath__63__W1[21]));
ADDHX1 cynw_cm_float_rcp_I2226 (.CO(N7410), .S(N7902), .A(inst_cellmath__62__W0[21]), .B(inst_cellmath__62__W1[21]));
ADDFX1 cynw_cm_float_rcp_I2227 (.CO(N7686), .S(N7552), .A(inst_cellmath__63__W0[22]), .B(N484), .CI(inst_cellmath__62__W0[22]));
ADDHX1 cynw_cm_float_rcp_I2228 (.CO(N7957), .S(N7817), .A(inst_cellmath__63__W1[22]), .B(inst_cellmath__62__W1[22]));
ADDFX1 cynw_cm_float_rcp_I2229 (.CO(N7606), .S(N7471), .A(inst_cellmath__62__W0[23]), .B(N485), .CI(inst_cellmath__62__W1[23]));
ADDHX1 cynw_cm_float_rcp_I2230 (.CO(N7874), .S(N7741), .A(inst_cellmath__63__W0[23]), .B(inst_cellmath__63__W1[23]));
ADDFX1 cynw_cm_float_rcp_I2231 (.CO(N7530), .S(N8010), .A(inst_cellmath__62__W0[24]), .B(N486), .CI(inst_cellmath__62__W1[24]));
ADDHX1 cynw_cm_float_rcp_I2232 (.CO(N7795), .S(N7659), .A(inst_cellmath__63__W0[24]), .B(inst_cellmath__63__W1[24]));
ADDHX1 cynw_cm_float_rcp_I2234 (.CO(N7719), .S(N7585), .A(inst_cellmath__63__W0[25]), .B(inst_cellmath__63__W1[25]));
ADDHX1 cynw_cm_float_rcp_I2236 (.CO(N7634), .S(N7508), .A(inst_cellmath__63__W0[26]), .B(inst_cellmath__63__W1[26]));
ADDHX1 cynw_cm_float_rcp_I2238 (.CO(N7563), .S(N7420), .A(inst_cellmath__63__W0[27]), .B(inst_cellmath__63__W1[27]));
ADDHX1 cynw_cm_float_rcp_I2240 (.CO(N7484), .S(N7965), .A(inst_cellmath__63__W0[28]), .B(inst_cellmath__63__W1[28]));
ADDHX1 cynw_cm_float_rcp_I2242 (.CO(N8018), .S(N7888), .A(inst_cellmath__63__W0[29]), .B(inst_cellmath__63__W1[29]));
ADDHX1 cynw_cm_float_rcp_I2244 (.CO(N7941), .S(N7803), .A(inst_cellmath__63__W0[30]), .B(inst_cellmath__63__W1[30]));
ADDHX1 cynw_cm_float_rcp_I2246 (.CO(N7862), .S(N7725), .A(inst_cellmath__63__W0[31]), .B(inst_cellmath__63__W1[31]));
ADDHX1 cynw_cm_float_rcp_I2248 (.CO(N7784), .S(N7645), .A(inst_cellmath__63__W0[32]), .B(inst_cellmath__63__W1[32]));
ADDHX1 cynw_cm_float_rcp_I2250 (.CO(N7706), .S(N7571), .A(N495), .B(inst_cellmath__63__W1[33]));
NOR4X1 cynw_cm_float_rcp_I5079 (.Y(N7909), .A(N6570), .B(N6301), .C(N6533), .D(N6077));
ADDHX1 cynw_cm_float_rcp_I2267 (.CO(N7562), .S(N7417), .A(inst_cellmath__63__W1[2]), .B(inst_cellmath__63__W0[2]));
ADDHX1 cynw_cm_float_rcp_I2269 (.CO(N7963), .S(N7823), .A(inst_cellmath__63__W1[3]), .B(inst_cellmath__63__W0[3]));
ADDHX1 cynw_cm_float_rcp_I2270 (.CO(N7884), .S(N7745), .A(inst_cellmath__63__W0[4]), .B(inst_cellmath__62__W0[4]));
ADDHX1 cynw_cm_float_rcp_I2271 (.CO(N7748), .S(N7612), .A(inst_cellmath__63__W1[4]), .B(N7745));
ADDFX1 cynw_cm_float_rcp_I2272 (.CO(N7667), .S(N7640), .A(inst_cellmath__62__W1[5]), .B(inst_cellmath__63__W0[5]), .CI(inst_cellmath__62__W0[5]));
ADDFX1 cynw_cm_float_rcp_I2273 (.CO(N7535), .S(N8016), .A(N7884), .B(inst_cellmath__63__W1[5]), .CI(N7640));
ADDFX1 cynw_cm_float_rcp_I2274 (.CO(N7451), .S(N7542), .A(inst_cellmath__63__W0[6]), .B(inst_cellmath__62__W0[6]), .CI(inst_cellmath__62__W1[6]));
ADDFX1 cynw_cm_float_rcp_I2275 (.CO(N7939), .S(N7802), .A(N7667), .B(inst_cellmath__63__W1[6]), .CI(N7542));
ADDFX1 cynw_cm_float_rcp_I2276 (.CO(N7857), .S(N7437), .A(inst_cellmath__63__W0[7]), .B(inst_cellmath__62__W0[7]), .CI(inst_cellmath__63__W1[7]));
ADDFX1 cynw_cm_float_rcp_I2277 (.CO(N7724), .S(N7592), .A(N7451), .B(inst_cellmath__62__W1[7]), .CI(N7437));
ADDFX1 cynw_cm_float_rcp_I2278 (.CO(N7643), .S(N7960), .A(inst_cellmath__62__W0[8]), .B(inst_cellmath__63__W0[8]), .CI(inst_cellmath__63__W1[8]));
ADDFX1 cynw_cm_float_rcp_I2279 (.CO(N7514), .S(N7995), .A(N7857), .B(inst_cellmath__62__W1[8]), .CI(N7960));
ADDFX1 cynw_cm_float_rcp_I2280 (.CO(N7429), .S(N7851), .A(inst_cellmath__63__W1[9]), .B(inst_cellmath__63__W0[9]), .CI(inst_cellmath__62__W0[9]));
ADDFX1 cynw_cm_float_rcp_I2281 (.CO(N7919), .S(N7780), .A(inst_cellmath__62__W1[9]), .B(N7643), .CI(N7851));
ADDFX1 cynw_cm_float_rcp_I2282 (.CO(N7832), .S(N7753), .A(inst_cellmath__63__W1[10]), .B(inst_cellmath__63__W0[10]), .CI(inst_cellmath__62__W0[10]));
ADDFX1 cynw_cm_float_rcp_I2283 (.CO(N7703), .S(N7570), .A(N7429), .B(inst_cellmath__62__W1[10]), .CI(N7753));
ADDFX1 cynw_cm_float_rcp_I2284 (.CO(N7622), .S(N7648), .A(inst_cellmath__63__W1[11]), .B(inst_cellmath__63__W0[11]), .CI(inst_cellmath__62__W0[11]));
ADDFX1 cynw_cm_float_rcp_I2285 (.CO(N7491), .S(N7971), .A(N7832), .B(inst_cellmath__62__W1[11]), .CI(N7648));
ADDFX1 cynw_cm_float_rcp_I2286 (.CO(N8024), .S(N7550), .A(inst_cellmath__63__W1[12]), .B(inst_cellmath__63__W0[12]), .CI(inst_cellmath__62__W0[12]));
ADDFX1 cynw_cm_float_rcp_I2287 (.CO(N7895), .S(N7761), .A(N7550), .B(N7622), .CI(inst_cellmath__62__W1[12]));
ADDFX1 cynw_cm_float_rcp_I2288 (.CO(N7811), .S(N7442), .A(inst_cellmath__63__W1[13]), .B(inst_cellmath__63__W0[13]), .CI(inst_cellmath__62__W0[13]));
ADDFX1 cynw_cm_float_rcp_I2289 (.CO(N7679), .S(N7545), .A(N8024), .B(inst_cellmath__62__W1[13]), .CI(N7442));
ADDFX1 cynw_cm_float_rcp_I2290 (.CO(N7601), .S(N7964), .A(inst_cellmath__63__W1[14]), .B(inst_cellmath__63__W0[14]), .CI(inst_cellmath__62__W0[14]));
ADDFX1 cynw_cm_float_rcp_I2291 (.CO(N7464), .S(N7952), .A(N7811), .B(inst_cellmath__62__W1[14]), .CI(N7964));
ADDFX1 cynw_cm_float_rcp_I2292 (.CO(N8005), .S(N7861), .A(inst_cellmath__63__W1[15]), .B(N7487), .CI(inst_cellmath__62__W0[15]));
ADDFXL cynw_cm_float_rcp_I2293 (.CO(N7869), .S(N7733), .A(N7601), .B(inst_cellmath__62__W1[15]), .CI(N7861));
ADDFHXL cynw_cm_float_rcp_I2294 (.CO(N7791), .S(N7763), .A(N7757), .B(N7618), .CI(inst_cellmath__62__W1[16]));
ADDFHXL cynw_cm_float_rcp_I2295 (.CO(N7653), .S(N7524), .A(N7675), .B(N8005), .CI(N7763));
ADDFX1 cynw_cm_float_rcp_I2296 (.CO(N7578), .S(N7655), .A(N7945), .B(N7890), .CI(N7806));
ADDFX1 cynw_cm_float_rcp_I2297 (.CO(N7439), .S(N7927), .A(N7791), .B(N7597), .CI(N7655));
ADDFXL cynw_cm_float_rcp_I2298 (.CO(N7984), .S(N7561), .A(N7864), .B(N7457), .CI(N7520));
ADDFXL cynw_cm_float_rcp_I2299 (.CO(N7844), .S(N7712), .A(N7578), .B(N7730), .CI(N7561));
ADDFX1 cynw_cm_float_rcp_I2300 (.CO(N7771), .S(N7450), .A(N7787), .B(N8001), .CI(N7434));
ADDFX1 cynw_cm_float_rcp_I2301 (.CO(N7631), .S(N7501), .A(N7984), .B(N7649), .CI(N7450));
ADDFX1 cynw_cm_float_rcp_I2302 (.CO(N7557), .S(N7969), .A(N7709), .B(N7924), .CI(N7575));
ADDFX1 cynw_cm_float_rcp_I2303 (.CO(N7415), .S(N7906), .A(N7771), .B(N7980), .CI(N7969));
ADDFX1 cynw_cm_float_rcp_I2304 (.CO(N7961), .S(N7868), .A(N7627), .B(N7838), .CI(N7902));
ADDFX1 cynw_cm_float_rcp_I2305 (.CO(N7821), .S(N7690), .A(N7557), .B(N7497), .CI(N7868));
ADDFX1 cynw_cm_float_rcp_I2306 (.CO(N7744), .S(N7770), .A(N7817), .B(N7767), .CI(N7552));
ADDFX1 cynw_cm_float_rcp_I2307 (.CO(N7610), .S(N7476), .A(N7961), .B(N7410), .CI(N7770));
ADDFX1 cynw_cm_float_rcp_I2308 (.CO(N7533), .S(N7663), .A(N7471), .B(N7741), .CI(N7686));
ADDFX1 cynw_cm_float_rcp_I2309 (.CO(N8013), .S(N7880), .A(N7744), .B(N7957), .CI(N7663));
ADDFX1 cynw_cm_float_rcp_I2310 (.CO(N7937), .S(N7565), .A(N7659), .B(N8010), .CI(N7874));
ADDFX1 cynw_cm_float_rcp_I2311 (.CO(N7799), .S(N7664), .A(N7533), .B(N7606), .CI(N7565));
ADDFX1 cynw_cm_float_rcp_I2312 (.CO(N7722), .S(N7459), .A(N7530), .B(N487), .CI(N7795));
ADDFX1 cynw_cm_float_rcp_I2313 (.CO(N7589), .S(N7447), .A(N7937), .B(N7585), .CI(N7459));
ADDHX1 cynw_cm_float_rcp_I2314 (.CO(N7511), .S(N7982), .A(N488), .B(N7508));
ADDFX1 cynw_cm_float_rcp_I2315 (.CO(N7992), .S(N7853), .A(N7722), .B(N7719), .CI(N7982));
ADDHX1 cynw_cm_float_rcp_I2316 (.CO(N7917), .S(N7876), .A(N489), .B(N7420));
ADDFX1 cynw_cm_float_rcp_I2317 (.CO(N7778), .S(N7638), .A(N7511), .B(N7634), .CI(N7876));
ADDHX1 cynw_cm_float_rcp_I2318 (.CO(N7700), .S(N7776), .A(N490), .B(N7965));
ADDFX1 cynw_cm_float_rcp_I2319 (.CO(N7568), .S(N7425), .A(N7917), .B(N7563), .CI(N7776));
ADDHX1 cynw_cm_float_rcp_I2320 (.CO(N7489), .S(N7674), .A(N491), .B(N7888));
ADDFX1 cynw_cm_float_rcp_I2321 (.CO(N7968), .S(N7829), .A(N7700), .B(N7484), .CI(N7674));
ADDHX1 cynw_cm_float_rcp_I2322 (.CO(N7892), .S(N7572), .A(N492), .B(N7803));
ADDFX1 cynw_cm_float_rcp_I2323 (.CO(N7758), .S(N7620), .A(N7489), .B(N8018), .CI(N7572));
ADDHX1 cynw_cm_float_rcp_I2324 (.CO(N7677), .S(N7468), .A(N493), .B(N7725));
ADDFX1 cynw_cm_float_rcp_I2325 (.CO(N7543), .S(N8022), .A(N7892), .B(N7941), .CI(N7468));
ADDHX1 cynw_cm_float_rcp_I2326 (.CO(N7460), .S(N7988), .A(N494), .B(N7645));
ADDFX1 cynw_cm_float_rcp_I2327 (.CO(N7947), .S(N7809), .A(N7677), .B(N7862), .CI(N7988));
ADDHX1 cynw_cm_float_rcp_I2328 (.CO(N7866), .S(N7886), .A(inst_cellmath__63__W0[33]), .B(N7571));
ADDFX1 cynw_cm_float_rcp_I2329 (.CO(N7732), .S(N7599), .A(N7460), .B(N7784), .CI(N7886));
ADDHX1 cynw_cm_float_rcp_I2330 (.CO(N7651), .S(N7783), .A(1'B1), .B(N496));
ADDFX1 cynw_cm_float_rcp_I2331 (.CO(N7523), .S(N8003), .A(N7866), .B(N7706), .CI(N7783));
XNOR2X1 hap1_A_I5096 (.Y(N7789), .A(N497), .B(N7651));
OR2XL hap1_A_I5097 (.Y(N7926), .A(N497), .B(N7651));
INVXL hap1_A_I14176 (.Y(N7582), .A(N498));
OR2XL hap1_A_I5099 (.Y(N7841), .A(1'B0), .B(N498));
INVXL hap1_A_I14177 (.Y(N7478), .A(N499));
OR2XL hap1_A_I5101 (.Y(N7629), .A(1'B0), .B(N499));
ADDHX1 cynw_cm_float_rcp_I2337 (.CO(N7499), .S(N7983), .A(N7841), .B(N7478));
XNOR2X1 hap1_A_I5102 (.Y(N7769), .A(N500), .B(N7629));
OR2XL hap1_A_I5103 (.Y(N7904), .A(N500), .B(N7629));
OR2XL cynw_cm_float_rcp_I5065 (.Y(N7894), .A(N3896), .B(a_man[22]));
NOR2XL cynw_cm_float_rcp_I2347 (.Y(N8012), .A(N7562), .B(N7823));
NAND2XL cynw_cm_float_rcp_I2348 (.Y(N7532), .A(N7562), .B(N7823));
AND2XL cynw_cm_float_rcp_I2350 (.Y(N7797), .A(N7963), .B(N7612));
NOR2XL cynw_cm_float_rcp_I2351 (.Y(N7936), .A(N7748), .B(N8016));
NAND2XL cynw_cm_float_rcp_I2352 (.Y(N7444), .A(N7748), .B(N8016));
AND2XL cynw_cm_float_rcp_I2354 (.Y(N7721), .A(N7535), .B(N7802));
NOR2XL cynw_cm_float_rcp_I2355 (.Y(N7849), .A(N7939), .B(N7592));
NAND2XL cynw_cm_float_rcp_I2356 (.Y(N7991), .A(N7939), .B(N7592));
AND2XL cynw_cm_float_rcp_I2358 (.Y(N7635), .A(N7724), .B(N7995));
NOR2XL cynw_cm_float_rcp_I2359 (.Y(N7777), .A(N7514), .B(N7780));
NAND2XL cynw_cm_float_rcp_I2360 (.Y(N7916), .A(N7514), .B(N7780));
AND2XL cynw_cm_float_rcp_I2362 (.Y(N7564), .A(N7919), .B(N7570));
NOR2XL cynw_cm_float_rcp_I2363 (.Y(N7699), .A(N7703), .B(N7971));
NAND2XL cynw_cm_float_rcp_I2364 (.Y(N7826), .A(N7703), .B(N7971));
AND2XL cynw_cm_float_rcp_I2366 (.Y(N7486), .A(N7491), .B(N7761));
NOR2XL cynw_cm_float_rcp_I2367 (.Y(N7615), .A(N7895), .B(N7545));
NAND2XL cynw_cm_float_rcp_I2368 (.Y(N7754), .A(N7895), .B(N7545));
NAND2XL cynw_cm_float_rcp_I5080 (.Y(N7998), .A(N7909), .B(N7417));
AOI21XL cynw_cm_float_rcp_I2373 (.Y(N7837), .A0(N7532), .A1(N7998), .B0(N8012));
OAI22XL cynw_cm_float_rcp_I5067 (.Y(N7605), .A0(N7797), .A1(N7837), .B0(N7963), .B1(N7612));
AOI21XL cynw_cm_float_rcp_I2377 (.Y(N7989), .A0(N7444), .A1(N7605), .B0(N7936));
OAI22XL cynw_cm_float_rcp_I5068 (.Y(N7670), .A0(N7721), .A1(N7989), .B0(N7535), .B1(N7802));
AOI21XL cynw_cm_float_rcp_I2381 (.Y(N7973), .A0(N7991), .A1(N7670), .B0(N7849));
OAI22XL cynw_cm_float_rcp_I5069 (.Y(N7583), .A0(N7635), .A1(N7973), .B0(N7724), .B1(N7995));
AOI21XL cynw_cm_float_rcp_I2385 (.Y(N7800), .A0(N7916), .A1(N7583), .B0(N7777));
OAI22XL cynw_cm_float_rcp_I5070 (.Y(N7948), .A0(N7564), .A1(N7800), .B0(N7919), .B1(N7570));
AOI21XL cynw_cm_float_rcp_I2389 (.Y(N7474), .A0(N7826), .A1(N7948), .B0(N7699));
OAI22XL cynw_cm_float_rcp_I5071 (.Y(N7540), .A0(N7486), .A1(N7474), .B0(N7491), .B1(N7761));
AO21XL cynw_cm_float_rcp_I2420 (.Y(N7419), .A0(N7540), .A1(N7754), .B0(N7615));
XOR2XL cynw_cm_float_rcp_I2421 (.Y(N7824), .A(N7679), .B(N7952));
XOR2XL cynw_cm_float_rcp_I2422 (.Y(N7481), .A(N7464), .B(N7733));
XOR2XL cynw_cm_float_rcp_I2423 (.Y(N7750), .A(N7869), .B(N7524));
OR2XL cynw_cm_float_rcp_I2424 (.Y(N7488), .A(N7653), .B(N7927));
XOR2XL cynw_cm_float_rcp_I2425 (.Y(N8017), .A(N7653), .B(N7927));
OR2XL cynw_cm_float_rcp_I2426 (.Y(N7807), .A(N7439), .B(N7712));
XOR2XL cynw_cm_float_rcp_I2427 (.Y(N7668), .A(N7439), .B(N7712));
OR2XL cynw_cm_float_rcp_I2428 (.Y(N7521), .A(N7501), .B(N7844));
XOR2XL cynw_cm_float_rcp_I2429 (.Y(N7940), .A(N7501), .B(N7844));
OR2XL cynw_cm_float_rcp_I2430 (.Y(N7840), .A(N7906), .B(N7631));
XOR2XL cynw_cm_float_rcp_I2431 (.Y(N7593), .A(N7906), .B(N7631));
OR2XL cynw_cm_float_rcp_I2432 (.Y(N7553), .A(N7415), .B(N7690));
XOR2XL cynw_cm_float_rcp_I2433 (.Y(N7858), .A(N7415), .B(N7690));
OR2XL cynw_cm_float_rcp_I2434 (.Y(N7875), .A(N7476), .B(N7821));
XOR2XL cynw_cm_float_rcp_I2435 (.Y(N7515), .A(N7476), .B(N7821));
OR2XL cynw_cm_float_rcp_I2436 (.Y(N7586), .A(N7880), .B(N7610));
XOR2XL cynw_cm_float_rcp_I2437 (.Y(N7782), .A(N7880), .B(N7610));
OR2XL cynw_cm_float_rcp_I2438 (.Y(N7914), .A(N7664), .B(N8013));
XOR2XL cynw_cm_float_rcp_I2439 (.Y(N7430), .A(N7664), .B(N8013));
OR2XL cynw_cm_float_rcp_I2440 (.Y(N7614), .A(N7447), .B(N7799));
XOR2XL cynw_cm_float_rcp_I2441 (.Y(N7704), .A(N7447), .B(N7799));
OR2XL cynw_cm_float_rcp_I2442 (.Y(N7942), .A(N7853), .B(N7589));
XOR2XL cynw_cm_float_rcp_I2443 (.Y(N7972), .A(N7853), .B(N7589));
OR2XL cynw_cm_float_rcp_I2444 (.Y(N7646), .A(N7638), .B(N7992));
XOR2XL cynw_cm_float_rcp_I2445 (.Y(N7623), .A(N7638), .B(N7992));
OR2XL cynw_cm_float_rcp_I2446 (.Y(N7976), .A(N7425), .B(N7778));
XOR2XL cynw_cm_float_rcp_I2447 (.Y(N7896), .A(N7425), .B(N7778));
OR2XL cynw_cm_float_rcp_I2448 (.Y(N7683), .A(N7829), .B(N7568));
XOR2XL cynw_cm_float_rcp_I2449 (.Y(N7546), .A(N7829), .B(N7568));
OR2XL cynw_cm_float_rcp_I2450 (.Y(N8009), .A(N7620), .B(N7968));
XOR2XL cynw_cm_float_rcp_I2451 (.Y(N7813), .A(N7620), .B(N7968));
OR2XL cynw_cm_float_rcp_I2452 (.Y(N7716), .A(N8022), .B(N7758));
XOR2XL cynw_cm_float_rcp_I2453 (.Y(N7465), .A(N8022), .B(N7758));
OR2XL cynw_cm_float_rcp_I2454 (.Y(N7418), .A(N7809), .B(N7543));
XOR2XL cynw_cm_float_rcp_I2455 (.Y(N7735), .A(N7809), .B(N7543));
OR2XL cynw_cm_float_rcp_I2456 (.Y(N7749), .A(N7599), .B(N7947));
XOR2XL cynw_cm_float_rcp_I2457 (.Y(N8006), .A(N7599), .B(N7947));
OR2XL cynw_cm_float_rcp_I2458 (.Y(N7452), .A(N8003), .B(N7732));
XOR2XL cynw_cm_float_rcp_I2459 (.Y(N7654), .A(N8003), .B(N7732));
OR2XL cynw_cm_float_rcp_I2460 (.Y(N7781), .A(N7789), .B(N7523));
XOR2XL cynw_cm_float_rcp_I2461 (.Y(N7929), .A(N7789), .B(N7523));
OR2XL cynw_cm_float_rcp_I2462 (.Y(N7492), .A(N7926), .B(N7582));
XOR2XL cynw_cm_float_rcp_I2463 (.Y(N7580), .A(N7926), .B(N7582));
NOR2XL cynw_cm_float_rcp_I2466 (.Y(N7985), .A(N7769), .B(N7499));
XOR2XL cynw_cm_float_rcp_I2467 (.Y(N7503), .A(N7769), .B(N7499));
XNOR2X1 cynw_cm_float_rcp_I2468 (.Y(N7772), .A(N7894), .B(N7904));
OAI2BB2XL cynw_cm_float_rcp_I2469 (.Y(N7558), .A0N(N7824), .A1N(N7419), .B0(N7679), .B1(N7952));
OAI2BB2X1 cynw_cm_float_rcp_I2470 (.Y(N7747), .A0N(N7481), .A1N(N7558), .B0(N7464), .B1(N7733));
OAI2BB2X1 cynw_cm_float_rcp_I2471 (.Y(N7590), .A0N(N7750), .A1N(N7747), .B0(N7869), .B1(N7524));
OAI2BB1XL cynw_cm_float_rcp_I2472 (.Y(N7702), .A0N(N8017), .A1N(N7590), .B0(N7488));
OAI2BB1X1 cynw_cm_float_rcp_I2473 (.Y(N7462), .A0N(N7668), .A1N(N7702), .B0(N7807));
OAI2BB1XL cynw_cm_float_rcp_I2474 (.Y(N7500), .A0N(N7940), .A1N(N7462), .B0(N7521));
OAI2BB1XL cynw_cm_float_rcp_I2475 (.Y(N7798), .A0N(N7593), .A1N(N7500), .B0(N7840));
OAI2BB1XL cynw_cm_float_rcp_I2476 (.Y(N7756), .A0N(N7858), .A1N(N7798), .B0(N7553));
OAI2BB1XL cynw_cm_float_rcp_I2477 (.Y(N7979), .A0N(N7515), .A1N(N7756), .B0(N7875));
OAI2BB1XL cynw_cm_float_rcp_I2478 (.Y(N7847), .A0N(N7782), .A1N(N7979), .B0(N7586));
OAI2BB1XL cynw_cm_float_rcp_I2479 (.Y(N7996), .A0N(N7430), .A1N(N7847), .B0(N7914));
OAI2BB1XL cynw_cm_float_rcp_I2480 (.Y(N7794), .A0N(N7704), .A1N(N7996), .B0(N7614));
OAI2BB1XL cynw_cm_float_rcp_I2481 (.Y(N7856), .A0N(N7972), .A1N(N7794), .B0(N7942));
OAI2BB1XL cynw_cm_float_rcp_I2482 (.Y(N7579), .A0N(N7623), .A1N(N7856), .B0(N7646));
OAI2BB1XL cynw_cm_float_rcp_I2483 (.Y(N7567), .A0N(N7896), .A1N(N7579), .B0(N7976));
OAI2BB1XL cynw_cm_float_rcp_I2484 (.Y(N7820), .A0N(N7546), .A1N(N7567), .B0(N7683));
OAI2BB1XL cynw_cm_float_rcp_I2485 (.Y(N7728), .A0N(N7813), .A1N(N7820), .B0(N8009));
OAI2BB1XL cynw_cm_float_rcp_I2486 (.Y(N7911), .A0N(N7465), .A1N(N7728), .B0(N7716));
OAI2BB1XL cynw_cm_float_rcp_I2487 (.Y(N7736), .A0N(N7735), .A1N(N7911), .B0(N7418));
OAI2BB1XL cynw_cm_float_rcp_I2488 (.Y(N7831), .A0N(N8006), .A1N(N7736), .B0(N7749));
OAI2BB1X1 cynw_cm_float_rcp_I2489 (.Y(N7588), .A0N(N7654), .A1N(N7831), .B0(N7452));
OAI2BB1X1 cynw_cm_float_rcp_I2490 (.Y(N7608), .A0N(N7929), .A1N(N7588), .B0(N7781));
OAI2BB1X1 cynw_cm_float_rcp_I2491 (.Y(N7899), .A0N(N7580), .A1N(N7608), .B0(N7492));
NAND2BX1 cynw_cm_float_rcp_I2492 (.Y(N7834), .AN(N7899), .B(N7983));
AO21XL cynw_cm_float_rcp_I2493 (.Y(N7427), .A0(N7503), .A1(N7834), .B0(N7985));
XNOR2X1 cynw_cm_float_rcp_I2497 (.Y(inst_cellmath__64[17]), .A(N7590), .B(N8017));
XNOR2X1 cynw_cm_float_rcp_I2498 (.Y(inst_cellmath__64[18]), .A(N7702), .B(N7668));
XNOR2X1 cynw_cm_float_rcp_I2499 (.Y(inst_cellmath__64[19]), .A(N7462), .B(N7940));
XNOR2X1 cynw_cm_float_rcp_I2500 (.Y(inst_cellmath__64[20]), .A(N7500), .B(N7593));
XNOR2X1 cynw_cm_float_rcp_I2501 (.Y(inst_cellmath__64[21]), .A(N7798), .B(N7858));
XNOR2X1 cynw_cm_float_rcp_I2502 (.Y(inst_cellmath__64[22]), .A(N7756), .B(N7515));
XNOR2X1 cynw_cm_float_rcp_I2503 (.Y(inst_cellmath__64[23]), .A(N7979), .B(N7782));
XNOR2X1 cynw_cm_float_rcp_I2504 (.Y(inst_cellmath__64[24]), .A(N7847), .B(N7430));
XNOR2X1 cynw_cm_float_rcp_I2505 (.Y(inst_cellmath__64[25]), .A(N7996), .B(N7704));
XNOR2X1 cynw_cm_float_rcp_I2506 (.Y(inst_cellmath__64[26]), .A(N7794), .B(N7972));
XNOR2X1 cynw_cm_float_rcp_I2507 (.Y(inst_cellmath__64[27]), .A(N7856), .B(N7623));
XNOR2X1 cynw_cm_float_rcp_I2508 (.Y(inst_cellmath__64[28]), .A(N7579), .B(N7896));
XNOR2X1 cynw_cm_float_rcp_I2509 (.Y(inst_cellmath__64[29]), .A(N7567), .B(N7546));
XNOR2X1 cynw_cm_float_rcp_I2510 (.Y(inst_cellmath__64[30]), .A(N7820), .B(N7813));
XNOR2X1 cynw_cm_float_rcp_I2511 (.Y(inst_cellmath__64[31]), .A(N7728), .B(N7465));
XNOR2X1 cynw_cm_float_rcp_I2512 (.Y(inst_cellmath__64[32]), .A(N7911), .B(N7735));
XNOR2X1 cynw_cm_float_rcp_I2513 (.Y(inst_cellmath__64[33]), .A(N7736), .B(N8006));
XNOR2X1 cynw_cm_float_rcp_I2514 (.Y(inst_cellmath__64[34]), .A(N7831), .B(N7654));
XNOR2X1 cynw_cm_float_rcp_I2515 (.Y(inst_cellmath__64[35]), .A(N7588), .B(N7929));
XNOR2X1 cynw_cm_float_rcp_I2516 (.Y(inst_cellmath__64[36]), .A(N7608), .B(N7580));
XNOR2X1 cynw_cm_float_rcp_I2517 (.Y(inst_cellmath__64[37]), .A(N7899), .B(N7983));
XNOR2X1 cynw_cm_float_rcp_I2518 (.Y(inst_cellmath__64[38]), .A(N7834), .B(N7503));
INVXL xor2_A_I5104 (.Y(N11788), .A(N7427));
MXI2XL xor2_A_I5105 (.Y(inst_cellmath__64[39]), .A(N11788), .B(N7427), .S0(N7772));
MX2XL inst_cellmath__68_0_I2520 (.Y(x[0]), .A(inst_cellmath__29), .B(inst_cellmath__64[17]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2521 (.Y(x[1]), .A(inst_cellmath__29), .B(inst_cellmath__64[18]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2522 (.Y(x[2]), .A(inst_cellmath__29), .B(inst_cellmath__64[19]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2523 (.Y(x[3]), .A(inst_cellmath__29), .B(inst_cellmath__64[20]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2524 (.Y(x[4]), .A(inst_cellmath__29), .B(inst_cellmath__64[21]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2525 (.Y(x[5]), .A(inst_cellmath__29), .B(inst_cellmath__64[22]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2526 (.Y(x[6]), .A(inst_cellmath__29), .B(inst_cellmath__64[23]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2527 (.Y(x[7]), .A(inst_cellmath__29), .B(inst_cellmath__64[24]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2528 (.Y(x[8]), .A(inst_cellmath__29), .B(inst_cellmath__64[25]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2529 (.Y(x[9]), .A(inst_cellmath__29), .B(inst_cellmath__64[26]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2530 (.Y(x[10]), .A(inst_cellmath__29), .B(inst_cellmath__64[27]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2531 (.Y(x[11]), .A(inst_cellmath__29), .B(inst_cellmath__64[28]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2532 (.Y(x[12]), .A(inst_cellmath__29), .B(inst_cellmath__64[29]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2533 (.Y(x[13]), .A(inst_cellmath__29), .B(inst_cellmath__64[30]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2534 (.Y(x[14]), .A(inst_cellmath__29), .B(inst_cellmath__64[31]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2535 (.Y(x[15]), .A(inst_cellmath__29), .B(inst_cellmath__64[32]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2536 (.Y(x[16]), .A(inst_cellmath__29), .B(inst_cellmath__64[33]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2537 (.Y(x[17]), .A(inst_cellmath__29), .B(inst_cellmath__64[34]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2538 (.Y(x[18]), .A(inst_cellmath__29), .B(inst_cellmath__64[35]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2539 (.Y(x[19]), .A(inst_cellmath__29), .B(inst_cellmath__64[36]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2540 (.Y(x[20]), .A(inst_cellmath__29), .B(inst_cellmath__64[37]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2541 (.Y(x[21]), .A(inst_cellmath__29), .B(inst_cellmath__64[38]), .S0(inst_cellmath__67));
INVXL mx2_A_I5106 (.Y(N11795), .A(inst_cellmath__67));
AO22XL mx2_A_I5107 (.Y(x[22]), .A0(inst_cellmath__29), .A1(N11795), .B0(inst_cellmath__64[39]), .B1(inst_cellmath__67));
assign inst_cellmath__19[1] = 1'B1;
assign inst_cellmath__19[2] = 1'B1;
assign inst_cellmath__19[3] = 1'B1;
assign inst_cellmath__19[4] = 1'B1;
assign inst_cellmath__19[5] = 1'B1;
assign inst_cellmath__19[6] = 1'B1;
assign inst_cellmath__19[7] = 1'B1;
assign inst_cellmath__19[8] = 1'B1;
assign inst_cellmath__20[2] = 1'B0;
assign inst_cellmath__20[4] = 1'B0;
assign inst_cellmath__20[6] = 1'B0;
assign inst_cellmath__51[18] = 1'B1;
assign inst_cellmath__60[0] = a_man[3];
assign inst_cellmath__60[1] = 1'B0;
assign inst_cellmath__60[2] = 1'B0;
assign inst_cellmath__60[3] = 1'B0;
assign inst_cellmath__60[4] = 1'B0;
assign inst_cellmath__60[5] = 1'B0;
assign inst_cellmath__60[6] = 1'B0;
assign inst_cellmath__60[7] = 1'B0;
assign inst_cellmath__60[8] = 1'B0;
assign inst_cellmath__60[9] = 1'B0;
assign inst_cellmath__60[10] = 1'B0;
assign inst_cellmath__60[11] = 1'B0;
assign inst_cellmath__60[12] = 1'B0;
assign inst_cellmath__60[13] = 1'B0;
assign inst_cellmath__60[14] = 1'B0;
assign inst_cellmath__60[15] = 1'B0;
assign inst_cellmath__60[16] = 1'B0;
assign inst_cellmath__60[17] = 1'B0;
assign inst_cellmath__60[18] = 1'B0;
assign inst_cellmath__60[19] = 1'B0;
assign inst_cellmath__60[20] = 1'B0;
assign inst_cellmath__62__W0[0] = 1'B0;
assign inst_cellmath__62__W0[1] = 1'B0;
assign inst_cellmath__62__W0[2] = 1'B0;
assign inst_cellmath__62__W0[3] = 1'B0;
assign inst_cellmath__62__W0[25] = 1'B0;
assign inst_cellmath__62__W0[26] = 1'B0;
assign inst_cellmath__62__W0[27] = 1'B0;
assign inst_cellmath__62__W0[28] = 1'B0;
assign inst_cellmath__62__W0[29] = 1'B0;
assign inst_cellmath__62__W0[30] = 1'B0;
assign inst_cellmath__62__W0[31] = 1'B0;
assign inst_cellmath__62__W0[32] = 1'B0;
assign inst_cellmath__62__W0[33] = 1'B0;
assign inst_cellmath__62__W0[34] = 1'B0;
assign inst_cellmath__62__W0[35] = 1'B0;
assign inst_cellmath__62__W0[36] = 1'B0;
assign inst_cellmath__62__W0[37] = 1'B0;
assign inst_cellmath__62__W0[38] = 1'B0;
assign inst_cellmath__62__W0[39] = 1'B0;
assign inst_cellmath__62__W1[0] = 1'B0;
assign inst_cellmath__62__W1[1] = 1'B0;
assign inst_cellmath__62__W1[2] = 1'B0;
assign inst_cellmath__62__W1[3] = 1'B0;
assign inst_cellmath__62__W1[4] = 1'B0;
assign inst_cellmath__62__W1[25] = 1'B0;
assign inst_cellmath__62__W1[26] = 1'B0;
assign inst_cellmath__62__W1[27] = 1'B0;
assign inst_cellmath__62__W1[28] = 1'B0;
assign inst_cellmath__62__W1[29] = 1'B0;
assign inst_cellmath__62__W1[30] = 1'B0;
assign inst_cellmath__62__W1[31] = 1'B0;
assign inst_cellmath__62__W1[32] = 1'B0;
assign inst_cellmath__62__W1[33] = 1'B0;
assign inst_cellmath__62__W1[34] = 1'B0;
assign inst_cellmath__62__W1[35] = 1'B0;
assign inst_cellmath__62__W1[36] = 1'B0;
assign inst_cellmath__62__W1[37] = 1'B0;
assign inst_cellmath__62__W1[38] = 1'B0;
assign inst_cellmath__62__W1[39] = 1'B0;
assign inst_cellmath__63__W0[0] = 1'B0;
assign inst_cellmath__63__W0[1] = 1'B0;
assign inst_cellmath__63__W0[34] = 1'B1;
assign inst_cellmath__63__W0[35] = 1'B1;
assign inst_cellmath__63__W0[36] = 1'B1;
assign inst_cellmath__63__W0[37] = 1'B1;
assign inst_cellmath__63__W0[38] = 1'B1;
assign inst_cellmath__63__W0[39] = 1'B1;
assign inst_cellmath__63__W1[0] = 1'B0;
assign inst_cellmath__63__W1[1] = 1'B0;
assign inst_cellmath__63__W1[34] = 1'B0;
assign inst_cellmath__63__W1[35] = 1'B0;
assign inst_cellmath__63__W1[36] = 1'B0;
assign inst_cellmath__63__W1[37] = 1'B0;
assign inst_cellmath__63__W1[38] = 1'B0;
assign inst_cellmath__63__W1[39] = 1'B0;
assign inst_cellmath__64[0] = 1'B0;
assign inst_cellmath__64[1] = 1'B0;
assign inst_cellmath__64[2] = 1'B0;
assign inst_cellmath__64[3] = 1'B0;
assign inst_cellmath__64[4] = 1'B0;
assign inst_cellmath__64[5] = 1'B0;
assign inst_cellmath__64[6] = 1'B0;
assign inst_cellmath__64[7] = 1'B0;
assign inst_cellmath__64[8] = 1'B0;
assign inst_cellmath__64[9] = 1'B0;
assign inst_cellmath__64[10] = 1'B0;
assign inst_cellmath__64[11] = 1'B0;
assign inst_cellmath__64[12] = 1'B0;
assign inst_cellmath__64[13] = 1'B0;
assign inst_cellmath__64[14] = 1'B0;
assign inst_cellmath__64[15] = 1'B0;
assign inst_cellmath__64[16] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  ubX0TwrdqB0= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



