/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:40:51 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__53,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__71,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4726,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4750,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4762,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4765,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7112,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755;
wire N5123,N5130,N5137,N5144,N5151,N5158,N5165 
	,N5172,N5179,N5186,N5193,N5200,N5207,N5214,N5221 
	,N5228,N5235,N5242,N5249,N5256,N5263,N5270,N5334 
	,N5336,N5572,N5585,N5587,N5611,N5613,N5676,N5683 
	,N5690,N5697,N5704,N5711,N5718,N5725,N5732,N5739 
	,N5746,N5753,N5760,N5767,N5774,N5781,N5788,N5795 
	,N5802,N5809,N5816,N5823,N5912,N5917,N5928,N5937 
	,N5946,N5955,N5964,N5973,N5982,N5991,N6000,N6153 
	,N6166,N6168,N6277,N6282,N6313,N6343,N6353,N6367 
	,N6369,N6400,N6419,N6425,N6427,N6451,N6456,N6458 
	,N6466,N6468,N6473,N6480,N6482,N6489,N6491,N6498 
	,N6507,N6509,N6516,N6525,N6527,N6534,N6543,N6545 
	,N6561,N6563,N6570,N6579,N6581,N6595,N6597,N6619 
	,N6649,N6688,N6737,N6794,N6851,N6909,N6967,N7025 
	,N7083,N7141,N7643,N7753,N7767,N7769,N7796,N7902 
	,N8095,N8097,N8099,N8182,N8198,N8261,N8556,N8564 
	,N8572,N8580,N8588,N8596,N8604,N8618,N8648,N8654 
	,N8663,N8670,N8677,N8684,N8691,N8699,N8707,N8715 
	,N8723,N8731,N8739,N8745,N8747,N8753,N8755,N8769 
	,N8779,N8781,N8787,N8797,N8799,N8805,N8815,N8817 
	,N8823,N8833,N8835,N8845,N8847,N8853,N8855,N8865 
	,N8867,N8873,N8875,N8885,N8887,N8893,N8895,N8905 
	,N8907,N8913,N8915,N8925,N8927,N8933,N8935,N8945 
	,N8947,N8953,N8955,N8965,N8967,N8977,N8981,N8983 
	,N9431,N9859;
reg x_reg_L0_22__retimed_I4673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4673_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1];
	end
assign N9431 = x_reg_L0_22__retimed_I4673_QOUT;
reg x_reg_L1_10__retimed_I4471_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I4471_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454;
	end
assign N8983 = x_reg_L1_10__retimed_I4471_QOUT;
reg x_reg_L1_10__retimed_I4470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I4470_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10];
	end
assign N8981 = x_reg_L1_10__retimed_I4470_QOUT;
reg x_reg_L1_9__retimed_I4468_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I4468_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9];
	end
assign N8977 = x_reg_L1_9__retimed_I4468_QOUT;
reg x_reg_L0_0__retimed_I4463_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4463_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657;
	end
assign N8967 = x_reg_L0_0__retimed_I4463_QOUT;
reg x_reg_L0_0__retimed_I4462_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4462_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3];
	end
assign N8965 = x_reg_L0_0__retimed_I4462_QOUT;
reg x_reg_L0_0__retimed_I4458_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4458_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658;
	end
assign N8955 = x_reg_L0_0__retimed_I4458_QOUT;
reg x_reg_L0_0__retimed_I4457_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4457_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4];
	end
assign N8953 = x_reg_L0_0__retimed_I4457_QOUT;
reg x_reg_L0_0__retimed_I4455_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4455_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659;
	end
assign N8947 = x_reg_L0_0__retimed_I4455_QOUT;
reg x_reg_L0_0__retimed_I4454_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4454_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5];
	end
assign N8945 = x_reg_L0_0__retimed_I4454_QOUT;
reg x_reg_L0_0__retimed_I4450_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4450_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660;
	end
assign N8935 = x_reg_L0_0__retimed_I4450_QOUT;
reg x_reg_L0_0__retimed_I4449_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4449_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6];
	end
assign N8933 = x_reg_L0_0__retimed_I4449_QOUT;
reg x_reg_L0_0__retimed_I4447_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4447_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7];
	end
assign N8927 = x_reg_L0_0__retimed_I4447_QOUT;
reg x_reg_L0_0__retimed_I4446_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4446_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661;
	end
assign N8925 = x_reg_L0_0__retimed_I4446_QOUT;
reg x_reg_L0_0__retimed_I4442_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4442_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662;
	end
assign N8915 = x_reg_L0_0__retimed_I4442_QOUT;
reg x_reg_L0_0__retimed_I4441_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4441_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8];
	end
assign N8913 = x_reg_L0_0__retimed_I4441_QOUT;
reg x_reg_L0_0__retimed_I4439_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4439_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663;
	end
assign N8907 = x_reg_L0_0__retimed_I4439_QOUT;
reg x_reg_L0_0__retimed_I4438_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4438_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9];
	end
assign N8905 = x_reg_L0_0__retimed_I4438_QOUT;
reg x_reg_L0_0__retimed_I4434_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4434_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664;
	end
assign N8895 = x_reg_L0_0__retimed_I4434_QOUT;
reg x_reg_L0_0__retimed_I4433_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4433_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10];
	end
assign N8893 = x_reg_L0_0__retimed_I4433_QOUT;
reg x_reg_L0_0__retimed_I4431_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4431_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665;
	end
assign N8887 = x_reg_L0_0__retimed_I4431_QOUT;
reg x_reg_L0_0__retimed_I4430_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4430_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11];
	end
assign N8885 = x_reg_L0_0__retimed_I4430_QOUT;
reg x_reg_L0_0__retimed_I4426_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4426_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666;
	end
assign N8875 = x_reg_L0_0__retimed_I4426_QOUT;
reg x_reg_L0_0__retimed_I4425_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4425_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12];
	end
assign N8873 = x_reg_L0_0__retimed_I4425_QOUT;
reg x_reg_L0_0__retimed_I4423_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4423_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667;
	end
assign N8867 = x_reg_L0_0__retimed_I4423_QOUT;
reg x_reg_L0_0__retimed_I4422_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4422_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13];
	end
assign N8865 = x_reg_L0_0__retimed_I4422_QOUT;
reg x_reg_L0_0__retimed_I4418_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4418_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668;
	end
assign N8855 = x_reg_L0_0__retimed_I4418_QOUT;
reg x_reg_L0_0__retimed_I4417_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4417_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14];
	end
assign N8853 = x_reg_L0_0__retimed_I4417_QOUT;
reg x_reg_L0_0__retimed_I4415_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4415_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669;
	end
assign N8847 = x_reg_L0_0__retimed_I4415_QOUT;
reg x_reg_L0_0__retimed_I4414_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4414_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15];
	end
assign N8845 = x_reg_L0_0__retimed_I4414_QOUT;
reg x_reg_L0_0__retimed_I4410_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4410_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670;
	end
assign N8835 = x_reg_L0_0__retimed_I4410_QOUT;
reg x_reg_L0_0__retimed_I4409_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4409_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16];
	end
assign N8833 = x_reg_L0_0__retimed_I4409_QOUT;
reg x_reg_L0_0__retimed_I4405_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4405_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588;
	end
assign N8823 = x_reg_L0_0__retimed_I4405_QOUT;
reg x_reg_L0_0__retimed_I4403_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4403_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672;
	end
assign N8817 = x_reg_L0_0__retimed_I4403_QOUT;
reg x_reg_L0_0__retimed_I4402_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4402_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18];
	end
assign N8815 = x_reg_L0_0__retimed_I4402_QOUT;
reg x_reg_L0_0__retimed_I4398_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4398_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568;
	end
assign N8805 = x_reg_L0_0__retimed_I4398_QOUT;
reg x_reg_L0_0__retimed_I4396_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4396_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674;
	end
assign N8799 = x_reg_L0_0__retimed_I4396_QOUT;
reg x_reg_L0_0__retimed_I4395_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4395_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20];
	end
assign N8797 = x_reg_L0_0__retimed_I4395_QOUT;
reg x_reg_L0_0__retimed_I4391_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4391_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550;
	end
assign N8787 = x_reg_L0_0__retimed_I4391_QOUT;
reg x_reg_L0_0__retimed_I4389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4389_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676;
	end
assign N8781 = x_reg_L0_0__retimed_I4389_QOUT;
reg x_reg_L0_0__retimed_I4388_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4388_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22];
	end
assign N8779 = x_reg_L0_0__retimed_I4388_QOUT;
reg x_reg_L0_0__retimed_I4384_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4384_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533;
	end
assign N8769 = x_reg_L0_0__retimed_I4384_QOUT;
reg x_reg_L0_0__retimed_I4379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4379_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541;
	end
assign N8755 = x_reg_L0_0__retimed_I4379_QOUT;
reg x_reg_L0_0__retimed_I4378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4378_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575;
	end
assign N8753 = x_reg_L0_0__retimed_I4378_QOUT;
reg x_reg_L0_0__retimed_I4377_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4377_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601;
	end
assign N8747 = x_reg_L0_0__retimed_I4377_QOUT;
reg x_reg_L0_0__retimed_I4376_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4376_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540;
	end
assign N8745 = x_reg_L0_0__retimed_I4376_QOUT;
reg x_reg_L0_0__retimed_I4375_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4375_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524;
	end
assign N8739 = x_reg_L0_0__retimed_I4375_QOUT;
reg x_reg_L0_0__retimed_I4373_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4373_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582;
	end
assign N8731 = x_reg_L0_0__retimed_I4373_QOUT;
reg x_reg_L0_0__retimed_I4371_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4371_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511;
	end
assign N8723 = x_reg_L0_0__retimed_I4371_QOUT;
reg x_reg_L0_0__retimed_I4369_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4369_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566;
	end
assign N8715 = x_reg_L0_0__retimed_I4369_QOUT;
reg x_reg_L0_0__retimed_I4367_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4367_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623;
	end
assign N8707 = x_reg_L0_0__retimed_I4367_QOUT;
reg x_reg_L0_0__retimed_I4365_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4365_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546;
	end
assign N8699 = x_reg_L0_0__retimed_I4365_QOUT;
reg x_reg_L0_0__retimed_I4363_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4363_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539;
	end
assign N8691 = x_reg_L0_0__retimed_I4363_QOUT;
reg x_reg_L0_0__retimed_I4361_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4361_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599;
	end
assign N8684 = x_reg_L0_0__retimed_I4361_QOUT;
reg x_reg_L0_0__retimed_I4359_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4359_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521;
	end
assign N8677 = x_reg_L0_0__retimed_I4359_QOUT;
reg x_reg_L0_0__retimed_I4357_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4357_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581;
	end
assign N8670 = x_reg_L0_0__retimed_I4357_QOUT;
reg x_reg_L0_0__retimed_I4355_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4355_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508;
	end
assign N8663 = x_reg_L0_0__retimed_I4355_QOUT;
reg x_reg_L0_0__retimed_I4352_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4352_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24];
	end
assign N8654 = x_reg_L0_0__retimed_I4352_QOUT;
reg x_reg_L0_0__retimed_I4351_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4351_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562;
	end
assign N8648 = x_reg_L0_0__retimed_I4351_QOUT;
reg x_reg_L0_0__retimed_I4342_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4342_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609;
	end
assign N8618 = x_reg_L0_0__retimed_I4342_QOUT;
reg x_reg_L0_0__retimed_I4338_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4338_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530;
	end
assign N8604 = x_reg_L0_0__retimed_I4338_QOUT;
reg x_reg_L0_0__retimed_I4336_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4336_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594;
	end
assign N8596 = x_reg_L0_0__retimed_I4336_QOUT;
reg x_reg_L0_0__retimed_I4334_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4334_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518;
	end
assign N8588 = x_reg_L0_0__retimed_I4334_QOUT;
reg x_reg_L0_0__retimed_I4332_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4332_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572;
	end
assign N8580 = x_reg_L0_0__retimed_I4332_QOUT;
reg x_reg_L0_0__retimed_I4330_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4330_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630;
	end
assign N8572 = x_reg_L0_0__retimed_I4330_QOUT;
reg x_reg_L0_0__retimed_I4328_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4328_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554;
	end
assign N8564 = x_reg_L0_0__retimed_I4328_QOUT;
reg x_reg_L0_0__retimed_I4326_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4326_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614;
	end
assign N8556 = x_reg_L0_0__retimed_I4326_QOUT;
reg x_reg_L0_0__retimed_I4222_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4222_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736;
	end
assign N8261 = x_reg_L0_0__retimed_I4222_QOUT;
reg x_reg_L0_0__retimed_I4197_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4197_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0];
	end
assign N8198 = x_reg_L0_0__retimed_I4197_QOUT;
reg x_reg_L0_0__retimed_I4192_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4192_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1];
	end
assign N8182 = x_reg_L0_0__retimed_I4192_QOUT;
reg x_reg_L0_0__retimed_I4173_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4173_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630;
	end
assign N8099 = x_reg_L0_0__retimed_I4173_QOUT;
reg x_reg_L0_0__retimed_I4172_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4172_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24];
	end
assign N8097 = x_reg_L0_0__retimed_I4172_QOUT;
reg x_reg_L0_0__retimed_I4171_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4171_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25];
	end
assign N8095 = x_reg_L0_0__retimed_I4171_QOUT;
reg x_reg_L0_0__retimed_I4136_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4136_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42;
	end
assign N7902 = x_reg_L0_0__retimed_I4136_QOUT;
reg x_reg_L0_0__retimed_I4112_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4112_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4;
	end
assign N7796 = x_reg_L0_0__retimed_I4112_QOUT;
reg x_reg_L0_0__retimed_I4102_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4102_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635;
	end
assign N7769 = x_reg_L0_0__retimed_I4102_QOUT;
reg x_reg_L0_0__retimed_I4101_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4101_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634;
	end
assign N7767 = x_reg_L0_0__retimed_I4101_QOUT;
reg x_reg_L0_0__retimed_I4095_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I4095_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557;
	end
assign N7753 = x_reg_L0_0__retimed_I4095_QOUT;
reg x_reg_L1_11__retimed_I4061_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I4061_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13];
	end
assign N7643 = x_reg_L1_11__retimed_I4061_QOUT;
reg x_reg_L1_12__retimed_I3866_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3866_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14];
	end
assign N7141 = x_reg_L1_12__retimed_I3866_QOUT;
reg x_reg_L1_13__retimed_I3843_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3843_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15];
	end
assign N7083 = x_reg_L1_13__retimed_I3843_QOUT;
reg x_reg_L1_14__retimed_I3820_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I3820_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16];
	end
assign N7025 = x_reg_L1_14__retimed_I3820_QOUT;
reg x_reg_L1_15__retimed_I3797_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3797_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17];
	end
assign N6967 = x_reg_L1_15__retimed_I3797_QOUT;
reg x_reg_L1_16__retimed_I3774_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3774_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18];
	end
assign N6909 = x_reg_L1_16__retimed_I3774_QOUT;
reg x_reg_L1_17__retimed_I3751_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3751_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19];
	end
assign N6851 = x_reg_L1_17__retimed_I3751_QOUT;
reg x_reg_L1_18__retimed_I3728_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3728_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20];
	end
assign N6794 = x_reg_L1_18__retimed_I3728_QOUT;
reg x_reg_L1_19__retimed_I3705_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3705_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21];
	end
assign N6737 = x_reg_L1_19__retimed_I3705_QOUT;
reg x_reg_L1_20__retimed_I3685_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I3685_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22];
	end
assign N6688 = x_reg_L1_20__retimed_I3685_QOUT;
reg x_reg_L1_21__retimed_I3669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I3669_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23];
	end
assign N6649 = x_reg_L1_21__retimed_I3669_QOUT;
reg x_reg_L1_22__retimed_I3657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I3657_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24];
	end
assign N6619 = x_reg_L1_22__retimed_I3657_QOUT;
reg x_reg_L1_23__retimed_I3649_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3649_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135;
	end
assign N6597 = x_reg_L1_23__retimed_I3649_QOUT;
reg x_reg_L1_23__retimed_I3648_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3648_QOUT <= N6570;
	end
assign N6595 = x_reg_L1_23__retimed_I3648_QOUT;
reg x_reg_L1_24__retimed_I3644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I3644_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614;
	end
assign N6581 = x_reg_L1_24__retimed_I3644_QOUT;
reg x_reg_L1_24__retimed_I3643_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I3643_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023;
	end
assign N6579 = x_reg_L1_24__retimed_I3643_QOUT;
reg x_reg_L0_22__retimed_I3640_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3640_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0];
	end
assign N6570 = x_reg_L0_22__retimed_I3640_QOUT;
reg x_reg_L1_25__retimed_I3638_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I3638_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079;
	end
assign N6563 = x_reg_L1_25__retimed_I3638_QOUT;
reg x_reg_L1_25__retimed_I3637_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I3637_QOUT <= N6534;
	end
assign N6561 = x_reg_L1_25__retimed_I3637_QOUT;
reg x_reg_L1_26__retimed_I3632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I3632_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158;
	end
assign N6545 = x_reg_L1_26__retimed_I3632_QOUT;
reg x_reg_L1_26__retimed_I3631_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I3631_QOUT <= N6516;
	end
assign N6543 = x_reg_L1_26__retimed_I3631_QOUT;
reg x_reg_L0_22__retimed_I3628_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3628_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605;
	end
assign N6534 = x_reg_L0_22__retimed_I3628_QOUT;
reg x_reg_L1_27__retimed_I3626_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I3626_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030;
	end
assign N6527 = x_reg_L1_27__retimed_I3626_QOUT;
reg x_reg_L1_27__retimed_I3625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I3625_QOUT <= N6498;
	end
assign N6525 = x_reg_L1_27__retimed_I3625_QOUT;
reg x_reg_L0_22__retimed_I3622_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3622_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630;
	end
assign N6516 = x_reg_L0_22__retimed_I3622_QOUT;
reg x_reg_L1_28__retimed_I3620_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I3620_QOUT <= N6482;
	end
assign N6509 = x_reg_L1_28__retimed_I3620_QOUT;
reg x_reg_L1_28__retimed_I3619_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I3619_QOUT <= N6480;
	end
assign N6507 = x_reg_L1_28__retimed_I3619_QOUT;
reg x_reg_L0_22__retimed_I3616_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3616_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600;
	end
assign N6498 = x_reg_L0_22__retimed_I3616_QOUT;
reg x_reg_L1_29__retimed_I3614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I3614_QOUT <= N6458;
	end
assign N6491 = x_reg_L1_29__retimed_I3614_QOUT;
reg x_reg_L1_29__retimed_I3613_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I3613_QOUT <= N6456;
	end
assign N6489 = x_reg_L1_29__retimed_I3613_QOUT;
reg x_reg_L0_22__retimed_I3611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3611_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612;
	end
assign N6482 = x_reg_L0_22__retimed_I3611_QOUT;
reg x_reg_L0_22__retimed_I3610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3610_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622;
	end
assign N6480 = x_reg_L0_22__retimed_I3610_QOUT;
reg x_reg_L1_12__retimed_I3608_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3608_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24];
	end
assign N6473 = x_reg_L1_12__retimed_I3608_QOUT;
reg x_reg_L1_30__retimed_I3606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I3606_QOUT <= N6427;
	end
assign N6468 = x_reg_L1_30__retimed_I3606_QOUT;
reg x_reg_L1_30__retimed_I3605_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I3605_QOUT <= N6425;
	end
assign N6466 = x_reg_L1_30__retimed_I3605_QOUT;
reg x_reg_L0_22__retimed_I3603_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3603_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617;
	end
assign N6458 = x_reg_L0_22__retimed_I3603_QOUT;
reg x_reg_L0_22__retimed_I3602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3602_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5];
	end
assign N6456 = x_reg_L0_22__retimed_I3602_QOUT;
reg x_reg_L1_12__retimed_I3601_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3601_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25];
	end
assign N6451 = x_reg_L1_12__retimed_I3601_QOUT;
reg x_reg_L0_22__retimed_I3591_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3591_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610;
	end
assign N6427 = x_reg_L0_22__retimed_I3591_QOUT;
reg x_reg_L0_22__retimed_I3590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3590_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6];
	end
assign N6425 = x_reg_L0_22__retimed_I3590_QOUT;
reg x_reg_L1_12__retimed_I3589_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3589_QOUT <= N6353;
	end
assign N6419 = x_reg_L1_12__retimed_I3589_QOUT;
reg x_reg_L1_12__retimed_I3582_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3582_QOUT <= N6343;
	end
assign N6400 = x_reg_L1_12__retimed_I3582_QOUT;
reg x_reg_L1_12__retimed_I3569_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3569_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5];
	end
assign N6369 = x_reg_L1_12__retimed_I3569_QOUT;
reg x_reg_L1_12__retimed_I3568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3568_QOUT <= N6313;
	end
assign N6367 = x_reg_L1_12__retimed_I3568_QOUT;
reg x_reg_L0_22__retimed_I3563_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3563_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134;
	end
assign N6353 = x_reg_L0_22__retimed_I3563_QOUT;
reg x_reg_L0_22__retimed_I3560_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3560_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7];
	end
assign N6343 = x_reg_L0_22__retimed_I3560_QOUT;
reg x_reg_L0_22__retimed_I3547_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3547_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189;
	end
assign N6313 = x_reg_L0_22__retimed_I3547_QOUT;
reg x_reg_L1_23__retimed_I3538_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3538_QOUT <= N5917;
	end
assign N6282 = x_reg_L1_23__retimed_I3538_QOUT;
reg x_reg_L1_22__retimed_I3536_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I3536_QOUT <= N5912;
	end
assign N6277 = x_reg_L1_22__retimed_I3536_QOUT;
reg x_reg_L1_23__retimed_I3522_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3522_QOUT <= N5587;
	end
assign N6168 = x_reg_L1_23__retimed_I3522_QOUT;
reg x_reg_L1_23__retimed_I3521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3521_QOUT <= N5585;
	end
assign N6166 = x_reg_L1_23__retimed_I3521_QOUT;
reg x_reg_L1_22__retimed_I3519_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I3519_QOUT <= N5572;
	end
assign N6153 = x_reg_L1_22__retimed_I3519_QOUT;
reg x_reg_L1_8__retimed_I3461_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3461_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8];
	end
assign N6000 = x_reg_L1_8__retimed_I3461_QOUT;
reg x_reg_L1_7__retimed_I3457_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3457_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7];
	end
assign N5991 = x_reg_L1_7__retimed_I3457_QOUT;
reg x_reg_L1_6__retimed_I3453_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3453_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6];
	end
assign N5982 = x_reg_L1_6__retimed_I3453_QOUT;
reg x_reg_L1_5__retimed_I3449_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3449_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5];
	end
assign N5973 = x_reg_L1_5__retimed_I3449_QOUT;
reg x_reg_L1_4__retimed_I3445_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3445_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4];
	end
assign N5964 = x_reg_L1_4__retimed_I3445_QOUT;
reg x_reg_L1_3__retimed_I3441_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3441_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3];
	end
assign N5955 = x_reg_L1_3__retimed_I3441_QOUT;
reg x_reg_L1_2__retimed_I3437_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3437_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2];
	end
assign N5946 = x_reg_L1_2__retimed_I3437_QOUT;
reg x_reg_L1_1__retimed_I3433_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3433_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1];
	end
assign N5937 = x_reg_L1_1__retimed_I3433_QOUT;
reg x_reg_L1_0__retimed_I3429_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3429_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0];
	end
assign N5928 = x_reg_L1_0__retimed_I3429_QOUT;
reg x_reg_L0_23__retimed_I3424_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3424_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650;
	end
assign N5917 = x_reg_L0_23__retimed_I3424_QOUT;
reg x_reg_L0_7__retimed_I3422_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I3422_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790;
	end
assign N5912 = x_reg_L0_7__retimed_I3422_QOUT;
reg x_reg_L1_0__retimed_I3413_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3413_QOUT <= N5270;
	end
assign N5823 = x_reg_L1_0__retimed_I3413_QOUT;
reg x_reg_L1_1__retimed_I3410_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3410_QOUT <= N5263;
	end
assign N5816 = x_reg_L1_1__retimed_I3410_QOUT;
reg x_reg_L1_2__retimed_I3407_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3407_QOUT <= N5256;
	end
assign N5809 = x_reg_L1_2__retimed_I3407_QOUT;
reg x_reg_L1_3__retimed_I3404_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3404_QOUT <= N5249;
	end
assign N5802 = x_reg_L1_3__retimed_I3404_QOUT;
reg x_reg_L1_4__retimed_I3401_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3401_QOUT <= N5242;
	end
assign N5795 = x_reg_L1_4__retimed_I3401_QOUT;
reg x_reg_L1_5__retimed_I3398_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3398_QOUT <= N5235;
	end
assign N5788 = x_reg_L1_5__retimed_I3398_QOUT;
reg x_reg_L1_6__retimed_I3395_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3395_QOUT <= N5228;
	end
assign N5781 = x_reg_L1_6__retimed_I3395_QOUT;
reg x_reg_L1_7__retimed_I3392_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3392_QOUT <= N5221;
	end
assign N5774 = x_reg_L1_7__retimed_I3392_QOUT;
reg x_reg_L1_8__retimed_I3389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3389_QOUT <= N5214;
	end
assign N5767 = x_reg_L1_8__retimed_I3389_QOUT;
reg x_reg_L1_9__retimed_I3386_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I3386_QOUT <= N5207;
	end
assign N5760 = x_reg_L1_9__retimed_I3386_QOUT;
reg x_reg_L1_10__retimed_I3383_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I3383_QOUT <= N5200;
	end
assign N5753 = x_reg_L1_10__retimed_I3383_QOUT;
reg x_reg_L1_11__retimed_I3380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I3380_QOUT <= N5193;
	end
assign N5746 = x_reg_L1_11__retimed_I3380_QOUT;
reg x_reg_L1_12__retimed_I3377_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3377_QOUT <= N5186;
	end
assign N5739 = x_reg_L1_12__retimed_I3377_QOUT;
reg x_reg_L1_13__retimed_I3374_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3374_QOUT <= N5179;
	end
assign N5732 = x_reg_L1_13__retimed_I3374_QOUT;
reg x_reg_L1_14__retimed_I3371_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I3371_QOUT <= N5172;
	end
assign N5725 = x_reg_L1_14__retimed_I3371_QOUT;
reg x_reg_L1_15__retimed_I3368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3368_QOUT <= N5165;
	end
assign N5718 = x_reg_L1_15__retimed_I3368_QOUT;
reg x_reg_L1_16__retimed_I3365_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3365_QOUT <= N5158;
	end
assign N5711 = x_reg_L1_16__retimed_I3365_QOUT;
reg x_reg_L1_17__retimed_I3362_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3362_QOUT <= N5151;
	end
assign N5704 = x_reg_L1_17__retimed_I3362_QOUT;
reg x_reg_L1_18__retimed_I3359_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3359_QOUT <= N5144;
	end
assign N5697 = x_reg_L1_18__retimed_I3359_QOUT;
reg x_reg_L1_19__retimed_I3356_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3356_QOUT <= N5137;
	end
assign N5690 = x_reg_L1_19__retimed_I3356_QOUT;
reg x_reg_L1_20__retimed_I3353_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I3353_QOUT <= N5130;
	end
assign N5683 = x_reg_L1_20__retimed_I3353_QOUT;
reg x_reg_L1_21__retimed_I3350_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I3350_QOUT <= N5123;
	end
assign N5676 = x_reg_L1_21__retimed_I3350_QOUT;
reg x_reg_L0_31__retimed_I3323_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3323_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6;
	end
assign N5613 = x_reg_L0_31__retimed_I3323_QOUT;
reg x_reg_L0_31__retimed_I3322_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3322_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
	end
assign N5611 = x_reg_L0_31__retimed_I3322_QOUT;
reg x_reg_L0_23__retimed_I3314_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3314_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12;
	end
assign N5587 = x_reg_L0_23__retimed_I3314_QOUT;
reg x_reg_L0_23__retimed_I3313_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3313_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17;
	end
assign N5585 = x_reg_L0_23__retimed_I3313_QOUT;
reg x_reg_L0_22__retimed_I3311_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3311_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
	end
assign N5572 = x_reg_L0_22__retimed_I3311_QOUT;
reg x_reg_L0_31__retimed_I3216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3216_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001;
	end
assign N5336 = x_reg_L0_31__retimed_I3216_QOUT;
reg x_reg_L0_31__retimed_I3215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3215_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010;
	end
assign N5334 = x_reg_L0_31__retimed_I3215_QOUT;
reg x_reg_L0_0__retimed_I3188_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I3188_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0];
	end
assign N5270 = x_reg_L0_0__retimed_I3188_QOUT;
reg x_reg_L0_1__retimed_I3185_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I3185_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1];
	end
assign N5263 = x_reg_L0_1__retimed_I3185_QOUT;
reg x_reg_L0_2__retimed_I3182_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I3182_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2];
	end
assign N5256 = x_reg_L0_2__retimed_I3182_QOUT;
reg x_reg_L0_3__retimed_I3179_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I3179_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3];
	end
assign N5249 = x_reg_L0_3__retimed_I3179_QOUT;
reg x_reg_L0_4__retimed_I3176_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I3176_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4];
	end
assign N5242 = x_reg_L0_4__retimed_I3176_QOUT;
reg x_reg_L0_5__retimed_I3173_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I3173_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5];
	end
assign N5235 = x_reg_L0_5__retimed_I3173_QOUT;
reg x_reg_L0_6__retimed_I3170_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I3170_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6];
	end
assign N5228 = x_reg_L0_6__retimed_I3170_QOUT;
reg x_reg_L0_7__retimed_I3167_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I3167_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7];
	end
assign N5221 = x_reg_L0_7__retimed_I3167_QOUT;
reg x_reg_L0_8__retimed_I3164_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I3164_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8];
	end
assign N5214 = x_reg_L0_8__retimed_I3164_QOUT;
reg x_reg_L0_9__retimed_I3161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I3161_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9];
	end
assign N5207 = x_reg_L0_9__retimed_I3161_QOUT;
reg x_reg_L0_10__retimed_I3158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I3158_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10];
	end
assign N5200 = x_reg_L0_10__retimed_I3158_QOUT;
reg x_reg_L0_11__retimed_I3155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I3155_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11];
	end
assign N5193 = x_reg_L0_11__retimed_I3155_QOUT;
reg x_reg_L0_12__retimed_I3152_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I3152_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12];
	end
assign N5186 = x_reg_L0_12__retimed_I3152_QOUT;
reg x_reg_L0_13__retimed_I3149_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I3149_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13];
	end
assign N5179 = x_reg_L0_13__retimed_I3149_QOUT;
reg x_reg_L0_14__retimed_I3146_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I3146_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14];
	end
assign N5172 = x_reg_L0_14__retimed_I3146_QOUT;
reg x_reg_L0_15__retimed_I3143_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I3143_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15];
	end
assign N5165 = x_reg_L0_15__retimed_I3143_QOUT;
reg x_reg_L0_16__retimed_I3140_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I3140_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16];
	end
assign N5158 = x_reg_L0_16__retimed_I3140_QOUT;
reg x_reg_L0_17__retimed_I3137_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I3137_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17];
	end
assign N5151 = x_reg_L0_17__retimed_I3137_QOUT;
reg x_reg_L0_18__retimed_I3134_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I3134_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18];
	end
assign N5144 = x_reg_L0_18__retimed_I3134_QOUT;
reg x_reg_L0_19__retimed_I3131_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I3131_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19];
	end
assign N5137 = x_reg_L0_19__retimed_I3131_QOUT;
reg x_reg_L0_20__retimed_I3128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I3128_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20];
	end
assign N5130 = x_reg_L0_20__retimed_I3128_QOUT;
reg x_reg_L0_21__retimed_I3125_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I3125_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21];
	end
assign N5123 = x_reg_L0_21__retimed_I3125_QOUT;
assign bdw_enable = !astall;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083 = !(a_exp[0] & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149 = !((a_exp[7] & a_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652 = !a_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653 | a_man[1]) | a_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106 = !(a_man[10] | a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125 = !(a_man[6] | a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114 = !(a_man[8] | a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134 = !(a_man[4] | a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168 = !(b_exp[0] & b_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157 = !((b_exp[7] & b_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208 = !(((b_man[0] | b_man[1]) | b_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191 = !(b_man[10] | b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210 = !(b_man[6] | b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199 = !(b_man[8] | b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219 = !(b_man[4] | b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25] = a_sign ^ b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563 = !b_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562 = !b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561 = !b_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560 = !b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559 = !b_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558 = !b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557 = !b_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556 = !b_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333 = a_exp[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1]} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2]} = {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3]} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4]} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5]} = {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6]} = {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7]} = {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7];
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556} + {1'B0, a_exp[0]};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364} + {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561} + {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562} + {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572} = {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638 = !a_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661 = b_man[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950 = !b_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633 = !(a_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642 = a_man[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459 = !a_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241 = !b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386 = !a_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387 = !b_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369 = !b_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371 = !a_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378 = !b_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384 = !a_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378 & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264 = !b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427 = !a_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428 = !b_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410 = !b_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412 = !a_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419 = !b_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425 = !a_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419 & a_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287 = !b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468 = !a_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469 = !b_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451 = !b_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453 = !a_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461 = !b_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466 = !a_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461 & a_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310 = !b_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319 = !a_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323 = !b_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346 = !a_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333 = !b_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351 = !b_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344 = !a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975 = !b_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975 | a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980 = !a_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985 = !(b_man[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986 = !a_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973 = !(b_man[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981 = !b_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977 = !(a_man[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980 & b_man[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323 & a_man[5]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314 & (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323 | a_man[5])));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319 & b_man[6]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317 & (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319 | b_man[6])));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310 & a_man[7]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321 & (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310 | a_man[7])));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466)) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430 = !((a_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298 & (a_man[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425)) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264 & a_man[15]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275 & (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264 | a_man[15])));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384)) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241 & a_man[19]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252 & (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241 | a_man[19])));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459 & b_man[20]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494 & (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459 | b_man[20])));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638 & b_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[20]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[19]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556 ^ a_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715 = !(N8182 | N8198);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510 = !((N8745 & N8747) | (!(N8965 | N8967)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592 = ((!N8739) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510)) | ((!N8953) & (!N8955));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592 & N8731) | (!(N8945 | N8947)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604 = ((!N8723) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537)) | ((!N8933) & (!N8935));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604 & N8715) | (!(N8925 | N8927)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585 = ((!N8707) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534)) | ((!N8913) & (!N8915));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585) ^ N8699;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534) ^ N8707;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604) ^ N8715;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537) ^ N8723;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592) ^ N8731;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510) ^ N8739;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3] = (!N8745) ^ N8747;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2] = (!N8753) ^ N8755;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585 & N8699) | (!(N8905 | N8907)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529 = ((!N8618) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631)) | ((!N8893) & (!N8895));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529 & N8604) | (!(N8885 | N8887)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576 = ((!N8596) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561)) | ((!N8873) & (!N8875));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576 & N8588) | (!(N8865 | N8867)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589 = ((!N8580) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593)) | ((!N8853) & (!N8855));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589 & N8572) | (!(N8845 | N8847)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564 = ((!N8564) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586)) | ((!N8833) & (!N8835));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564) ^ N8556;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586) ^ N8564;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589) ^ N8572;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593) ^ N8580;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576) ^ N8588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561) ^ N8596;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529) ^ N8604;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631) ^ N8618;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564 & N8556) | N8823);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512 = ((!N8691) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544)) | ((!N8815) & (!N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512 & N8684) | N8805);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549 = ((!N8677) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605)) | ((!N8797) & (!N8799));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549) ^ N8670;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605) ^ N8677;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512) ^ N8684;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544) ^ N8691;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549 & N8670) | N8787);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629) ^ N8663;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558 = ((!N8663) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629)) | ((!N8779) & (!N8781));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558) ^ N8648;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558 & N8648) | N8769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622) ^ N8654;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4617 = !(N8654 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7112 = N8095 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4617;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7112;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4750 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4750);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751 = !((N8261 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4762 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4790 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4765 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4762) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4790);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4726 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4754 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4805 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4726)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4754);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4793 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4765 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4805);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4793));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4716 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780;
assign N9859 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4716;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158 = (!N9859) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N8198);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102 = N8182 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031 = N8198 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N8182);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43 = (N8095 & N8099) | ((!N8095) & N8097);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__53 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582 | (!a_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565 = b_sign & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585 = !rm[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547 = !rm[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374 = !(N7902 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12550 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558) & N7902));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12592 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12560 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12550 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12592);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585 & rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5 = !(rm[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582 & b_sign) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582) & a_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12578 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12560 & N7796) | N7769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N636 = !(N7753 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12578);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__54 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558) & N7902);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N639 = ((!N7769) & (!N7767)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N639) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__53 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N636);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]} = {1'B0, N7643} + {1'B0, N8983};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]} = {1'B0, N7141} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]} = {1'B0, N7083} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]} = {1'B0, N7025} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]} = {1'B0, N6967} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]} = {1'B0, N6909} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]} = {1'B0, N6851} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]} = {1'B0, N6794} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]} = {1'B0, N6737} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]} = {1'B0, N6688} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]} = {1'B0, N6649} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23], fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]} = {1'B0, N6619} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151 = N6473 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151 | N6451);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755 | N6419);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6];
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614 = !N9431;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12123, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]} = {1'B0, N6595} + {1'B0, N6597} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12160, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]} = {1'B0, N6579} + {1'B0, N6581} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12123};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12194, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]} = {1'B0, N6561} + {1'B0, N6563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12160};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12148, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]} = {1'B0, N6543} + {1'B0, N6545} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12194};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12184, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]} = {1'B0, N6525} + {1'B0, N6527} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12148};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12139, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]} = {1'B0, N6507} + {1'B0, N6509} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12184};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12174, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]} = {1'B0, N6489} + {1'B0, N6491} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12139};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]} = {1'B0, N6466} + {1'B0, N6468} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12174};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12165 = !(N6400 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12125 = !(((N6367 | N6369) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12165);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12157 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12188 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12145 = (!N6400) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12177 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12188 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12145);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12162 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12157 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12177);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__71 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12125 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12162);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__71;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 | (!N6153));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769 = !(rm[0] & rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7 = !(rm[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70 = N6277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 = !(N6153 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]));
assign x[22] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[21]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]));
assign x[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5676);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[20]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]));
assign x[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5683);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[19]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]));
assign x[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5690);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[18]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]));
assign x[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5697);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[17]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]));
assign x[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5704);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[16]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]));
assign x[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5711);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[15]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]));
assign x[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[14]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]));
assign x[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5725);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[13]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]));
assign x[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5732);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[12]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]));
assign x[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5739);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[11]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]));
assign x[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5746);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[10]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & N8981));
assign x[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5753);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[9]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & N8977));
assign x[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5760);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[8]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & N6000));
assign x[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5767);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[7]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5991));
assign x[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5774);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[6]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5982));
assign x[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5781);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[5]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5973));
assign x[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5788);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[4]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5964));
assign x[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5795);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[3]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5955));
assign x[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5802);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5946));
assign x[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5809);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5937));
assign x[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5816);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & N5928));
assign x[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N5823);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745 = ((N6168 | N6166) | N6153) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751;
assign x[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]);
assign x[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]);
assign x[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]);
assign x[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]);
assign x[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]);
assign x[25] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]);
assign x[24] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651 = N6282 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0] = ((N6166 | N6168) | N6153) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651;
assign x[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748 = a_sign | b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6) | (a_sign & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_sign) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5] & N5613) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]) & N5611);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[31] = (N5334 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004) | ((!N5334) & N5336);
reg x_reg_L1_31__I1040_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I1040_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[31];
	end
assign x[31] = x_reg_L1_31__I1040_QOUT;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[0] = x[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[1] = x[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[2] = x[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[3] = x[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[4] = x[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[5] = x[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[6] = x[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[7] = x[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[8] = x[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[9] = x[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[10] = x[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[11] = x[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[12] = x[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[13] = x[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[14] = x[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[15] = x[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[16] = x[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[17] = x[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[18] = x[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[19] = x[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[20] = x[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[21] = x[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[22] = x[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[23] = x[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[24] = x[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[25] = x[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[26] = x[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[27] = x[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[28] = x[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[29] = x[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[30] = x[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[29] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[35] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[39] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  uLX3Sgncrxk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/


