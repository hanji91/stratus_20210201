/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:37:39 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_0_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__8,
	inst_cellmath__9,
	inst_cellmath__10,
	inst_cellmath__11,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__16,
	inst_cellmath__17,
	inst_cellmath__18;
wire [8:0] inst_cellmath__27;
wire [7:0] inst_cellmath__29;
wire  inst_cellmath__30;
wire [49:0] inst_cellmath__33;
wire [7:0] inst_cellmath__35;
wire [49:0] inst_cellmath__36,
	inst_cellmath__37;
wire [25:0] inst_cellmath__39;
wire  inst_cellmath__43,
	inst_cellmath__44;
wire [26:0] inst_cellmath__45;
wire  inst_cellmath__48;
wire [5:0] inst_cellmath__49;
wire [24:0] inst_cellmath__50;
wire  inst_cellmath__53,
	inst_cellmath__54,
	inst_cellmath__55;
wire [23:0] inst_cellmath__57;
wire [9:0] inst_cellmath__59;
wire  inst_cellmath__62,
	inst_cellmath__63;
wire [22:0] inst_cellmath__64;
wire  inst_cellmath__66;
wire [7:0] inst_cellmath__68;
wire  inst_cellmath__70,
	inst_cellmath__71;
wire N556,N557,N558,N559,N560,N561,N562 
	,N563,N565,N566,N567,N569,N570,N571,N572 
	,N573,N626,N627,N634,N635,N639,N642,N645 
	,N651,N652,N655,N656,N657,N658,N659,N660 
	,N661,N662,N663,N664,N665,N666,N667,N668 
	,N669,N671,N672,N673,N674,N675,N676,N677 
	,N706,N710,N1693,N2855,N4309,N4317,N4321,N4338 
	,N4340,N4346,N4352,N4354,N4357,N4369,N4373,N4377 
	,N4379,N4412,N4416,N4433,N4437,N4447,N4454,N4462 
	,N4464,N4468,N4474,N4525,N4581,N4582,N4591,N4592 
	,N4594,N4595,N4596,N4598,N4601,N4602,N4603,N4606 
	,N4607,N4609,N4610,N4611,N4613,N4614,N4615,N4617 
	,N4619,N4621,N4623,N4624,N4625,N4626,N4627,N4630 
	,N4631,N4634,N4635,N4637,N4638,N4640,N4641,N4643 
	,N4645,N4647,N4648,N4649,N4650,N4654,N4656,N4658 
	,N4659,N4661,N4662,N4664,N4665,N4666,N4667,N4668 
	,N4671,N4673,N4674,N4676,N4677,N4678,N4680,N4682 
	,N4684,N4685,N4687,N4688,N4690,N4692,N4695,N4697 
	,N4789,N4790,N4791,N4792,N4794,N4796,N4799,N4800 
	,N4801,N4802,N4805,N4806,N4807,N4809,N4810,N4812 
	,N4814,N4816,N4817,N4818,N4819,N4820,N4822,N4823 
	,N4824,N4825,N4828,N4829,N4830,N4832,N4835,N4836 
	,N4837,N4839,N4840,N4841,N4843,N4845,N4846,N4847 
	,N4848,N4851,N4853,N4854,N4856,N4857,N4859,N4861 
	,N4863,N4864,N4865,N4866,N4868,N4869,N4871,N4873 
	,N4874,N4875,N4876,N4878,N4880,N4881,N4882,N4884 
	,N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4897 
	,N4898,N4899,N4901,N4903,N4904,N4906,N4908,N4910 
	,N4911,N4912,N4914,N4915,N4917,N4919,N4921,N4922 
	,N4923,N4924,N4926,N4927,N4928,N4929,N4931,N4933 
	,N4934,N4935,N4938,N5094,N5114,N5119,N5123,N5141 
	,N5148,N5153,N5164,N5168,N5175,N5180,N5184,N5191 
	,N5195,N5201,N5206,N5210,N5217,N5222,N5224,N5233 
	,N5237,N5244,N5249,N5253,N5259,N5336,N5338,N5340 
	,N5342,N5345,N5346,N5347,N5348,N5350,N5352,N5355 
	,N5357,N5359,N5360,N5362,N5363,N5365,N5366,N5367 
	,N5372,N5373,N5375,N5376,N5377,N5379,N5382,N5383 
	,N5385,N5387,N5390,N5391,N5394,N5395,N5396,N5397 
	,N5398,N5401,N5405,N5406,N5407,N5409,N5412,N5415 
	,N5416,N5418,N5420,N5423,N5424,N5426,N5428,N5429 
	,N5431,N5434,N5436,N5438,N5440,N5441,N5443,N5445 
	,N5447,N5450,N5452,N5454,N5458,N5459,N5461,N5464 
	,N5467,N5468,N5470,N5471,N5473,N5474,N5479,N5480 
	,N5482,N5485,N5486,N5489,N5490,N5492,N5495,N5496 
	,N5498,N5499,N5501,N5503,N5504,N5505,N5506,N5511 
	,N5513,N5515,N5518,N5519,N5521,N5523,N5525,N5527 
	,N5529,N5531,N5534,N5535,N5536,N5538,N5541,N5544 
	,N5545,N5547,N5548,N5551,N5554,N5555,N5558,N5559 
	,N5560,N5562,N5563,N5567,N5568,N5569,N5571,N5574 
	,N5577,N5578,N5579,N5581,N5583,N5837,N5890,N5892 
	,N5894,N5899,N5901,N5905,N5909,N5916,N5919,N5922 
	,N5924,N5926,N5931,N5955,N5967,N6017,N6023,N6154 
	,N6155,N6156,N6158,N6159,N6160,N6161,N6162,N6164 
	,N6165,N6166,N6167,N6168,N6170,N6172,N6173,N6174 
	,N6176,N6177,N6178,N6179,N6180,N6182,N6184,N6185 
	,N6186,N6187,N6188,N6189,N6191,N6192,N6194,N6195 
	,N6197,N6198,N6199,N6200,N6201,N6202,N6204,N6205 
	,N6207,N6208,N6209,N6210,N6211,N6213,N6214,N6215 
	,N6217,N6218,N6220,N6222,N6223,N6225,N6226,N6227 
	,N6228,N6229,N6232,N6233,N6234,N6235,N6236,N6238 
	,N6239,N6240,N6242,N6244,N6245,N6247,N6248,N6249 
	,N6250,N6251,N6252,N6253,N6254,N6256,N6258,N6260 
	,N6261,N6262,N6263,N6264,N6266,N6267,N6268,N6270 
	,N6272,N6273,N6274,N6275,N6277,N6278,N6279,N6280 
	,N6281,N6282,N6284,N6286,N6287,N6288,N6291,N6292 
	,N6293,N6294,N6295,N6296,N6298,N6300,N6302,N6303 
	,N6304,N6305,N6307,N6308,N6310,N6311,N6312,N6314 
	,N6315,N6316,N6317,N6318,N6320,N6321,N6323,N6324 
	,N6325,N6327,N6328,N6329,N6330,N6331,N6334,N6335 
	,N6336,N6338,N6339,N6340,N6341,N6342,N6344,N6346 
	,N6347,N6348,N6349,N6350,N6351,N6352,N6353,N6354 
	,N6355,N6357,N6359,N6360,N6362,N6363,N6364,N6365 
	,N6366,N6367,N6369,N6371,N6372,N6373,N6374,N6375 
	,N6376,N6377,N6379,N6380,N6381,N6382,N6384,N6386 
	,N6387,N6388,N6390,N6391,N6392,N6393,N6394,N6395 
	,N6397,N6400,N6401,N6402,N6403,N6404,N6406,N6408 
	,N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6418 
	,N6419,N6421,N6422,N6423,N6424,N6426,N6428,N6429 
	,N6430,N6432,N6434,N6435,N6436,N6437,N6439,N6440 
	,N6441,N6442,N6443,N6446,N6447,N6448,N6449,N6450 
	,N6451,N6452,N6454,N6456,N6457,N6459,N6460,N6461 
	,N6462,N6463,N6464,N6465,N6466,N6467,N6469,N6471 
	,N6472,N6473,N6474,N6475,N6476,N6477,N6478,N6480 
	,N6760,N6762,N6763,N6764,N6765,N6768,N6769,N6772 
	,N6773,N6774,N6775,N6777,N6778,N6779,N6782,N6783 
	,N6785,N6787,N6790,N6793,N6794,N6795,N6797,N6798 
	,N6800,N6801,N6802,N6804,N6806,N6807,N6808,N6810 
	,N6811,N6812,N6815,N6816,N6818,N6819,N6821,N6823 
	,N6825,N6826,N6827,N6829,N6830,N6831,N6832,N6834 
	,N6836,N6838,N6839,N6840,N6842,N6843,N6845,N6847 
	,N6848,N6849,N6851,N6852,N6855,N6856,N6958,N6966 
	,N6969,N6977,N6984,N6987,N6995,N7000,N7004,N7011 
	,N7016,N7017,N7025,N7028,N7034,N7035,N7042,N7045 
	,N7050,N7054,N7060,N7064,N7071,N7076,N7086,N7090 
	,N7092,N7096,N7182,N7185,N7191,N7197,N7198,N7199 
	,N7200,N7202,N7204,N7206,N7207,N7208,N7209,N7211 
	,N7214,N7215,N7216,N7218,N7219,N7221,N7222,N7224 
	,N7225,N7228,N7229,N7230,N7232,N7234,N7235,N7236 
	,N7237,N7238,N7240,N7242,N7243,N7244,N7246,N7247 
	,N7251,N7252,N7253,N7255,N7257,N7258,N7260,N7261 
	,N7263,N7265,N7266,N7267,N7269,N7272,N7273,N7274 
	,N7276,N7277,N7279,N7280,N7282,N7284,N7286,N7287 
	,N7289,N7290,N7292,N7294,N7295,N7297,N7298,N7301 
	,N7303,N7304,N7305,N7308,N7310,N7312,N7313,N7315 
	,N7316,N7317,N7319,N7322,N7323,N7324,N7326,N7327 
	,N7329,N7330,N7331,N7333,N7335,N7336,N7339,N7340 
	,N7341,N7342,N7345,N7346,N7348,N7349,N7351,N7352 
	,N7354,N7357,N7359,N7360,N7361,N7363,N7503,N7524 
	,N7530,N7558,N7567,N7603,N7606,N7625,N7640,N7647 
	,N7661,N7667,N7668,N7670,N7671,N7672,N7675,N7676 
	,N7678,N7679,N7682,N7684,N7686,N7688,N7689,N7691 
	,N7693,N7694,N7695,N7696,N7699,N7701,N7702,N7704 
	,N7705,N7706,N7708,N7710,N7712,N7713,N7716,N7717 
	,N7718,N7721,N7722,N7724,N7728,N7729,N7731,N7732 
	,N7735,N7737,N7739,N7741,N7742,N7746,N7747,N7748 
	,N7751,N7753,N7754,N7755,N7757,N7758,N7759,N7761 
	,N7763,N7766,N7768,N7769,N7772,N7773,N7775,N7776 
	,N7781,N7782,N7786,N7788,N7791,N7792,N7795,N7796 
	,N7797,N7798,N7800,N7801,N7803,N7804,N7806,N7808 
	,N7941,N7945,N7946,N7950,N7961,N7970,N7972,N7976 
	,N7980,N8015,N8021,N8024,N8025,N8034,N8037,N8038 
	,N8042,N8044,N8045,N8048,N8049,N8053,N8055,N8056 
	,N8057,N8058,N8059,N8062,N8064,N8066,N8067,N8068 
	,N8070,N8071,N8072,N8074,N8075,N8076,N8078,N8079 
	,N8080,N8081,N8082,N8083,N8084,N8086,N8087,N8088 
	,N8090,N8094,N8099,N8100,N8101,N8104,N8106,N8107 
	,N8109,N8110,N8111,N8112,N8115,N8116,N8118,N8243 
	,N8253,N8276,N8296,N8317,N8339,N8346,N8353,N8358 
	,N8363,N8368,N8373,N8379,N8384,N8388,N8394,N8400 
	,N8407,N8412,N8417,N8424,N8426,N8429,N8435,N8440 
	,N8445,N8451,N8456,N8461,N8466,N10715,N10721,N10733 
	,N10734,N10735,N10736,N10737,N10738,N10742,N10745,N10761 
	,N10769,N10775,N10782,N10790,N10794,N10801,N10808,N10815 
	,N10822,N10829,N10836,N10843,N10851,N10862,N10869,N17371 
	,N17372,N17379,N17391,N17393,N17456,N17458,N17463,N17466 
	,N17470,N17475,N17480,N17483,N17485,N17489,N17493,N17513 
	,N17517,N17525,N17529,N17535,N17541,N17569,N17571,N17576 
	,N17578,N17580,N17583,N17586,N17588,N17590,N17592,N17595 
	,N17597,N17618,N17620,N17626,N17628,N17631,N17632,N17637 
	,N17638,N17642,N17644,N17648,N17649,N17653,N17655,N17660 
	,N17663,N17664,N17746,N17752,N17754,N17767,N17769,N17776 
	,N17778,N17805,N17808,N17811,N17814,N17818,N17821,N17825 
	,N17828,N17829,N17830,N17835,N17851,N17859,N17869,N17895 
	,N17922,N17933,N17945,N17952,N17959,N17966,N17974,N17979 
	;
AND4XL inst_cellmath__9_0_I11219 (.Y(N4317), .A(a_exp[0]), .B(a_exp[1]), .C(a_exp[7]), .D(a_exp[6]));
AND4XL inst_cellmath__9_0_I11220 (.Y(N4321), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND2XL inst_cellmath__9_0_I810 (.Y(inst_cellmath__9), .A(N4317), .B(N4321));
NOR2XL inst_cellmath__10__1__I812 (.Y(N4377), .A(a_man[22]), .B(a_man[21]));
NOR2XL inst_cellmath__10__1__I813 (.Y(N4340), .A(a_man[20]), .B(a_man[19]));
NOR2XL inst_cellmath__10__1__I819 (.Y(N4354), .A(a_man[8]), .B(a_man[7]));
INVX2 inst_cellmath__10__1__I822 (.Y(N4338), .A(a_man[2]));
OR4X1 inst_cellmath__10__1__I11221 (.Y(N4369), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__10__1__I11222 (.Y(N4379), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR2XL inst_cellmath__10__1__I830 (.Y(N4373), .A(N4369), .B(N4379));
NAND3XL hyperpropagate_4_1_A_I4737 (.Y(N10761), .A(N4377), .B(N4373), .C(N4340));
NOR4BX1 hyperpropagate_4_1_A_I11225 (.Y(N4346), .AN(N4338), .B(a_man[0]), .C(N10761), .D(a_man[1]));
OR4X1 inst_cellmath__10__1__I11224 (.Y(N4352), .A(a_man[6]), .B(a_man[4]), .C(a_man[5]), .D(a_man[3]));
NOR4BX1 inst_cellmath__10__1__I11226 (.Y(N4357), .AN(N4354), .B(a_man[10]), .C(N4352), .D(a_man[9]));
NAND2XL inst_cellmath__10__1__I833 (.Y(inst_cellmath__10), .A(N4357), .B(N4346));
NOR2XL cynw_cm_float_add2_ieee_I834 (.Y(inst_cellmath__12), .A(inst_cellmath__9), .B(inst_cellmath__10));
AND4XL inst_cellmath__14_0_I11227 (.Y(N4412), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[7]), .D(b_exp[6]));
AND4XL inst_cellmath__14_0_I11228 (.Y(N4416), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND2XL inst_cellmath__14_0_I841 (.Y(inst_cellmath__14), .A(N4412), .B(N4416));
NOR2XL inst_cellmath__15__3__I842 (.Y(N4462), .A(b_man[0]), .B(b_man[1]));
INVXL inst_cellmath__15__3__I853 (.Y(N4433), .A(b_man[2]));
OR4X1 inst_cellmath__15__3__I11229 (.Y(N4454), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__15__3__I11230 (.Y(N4464), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__15__3__I11231 (.Y(N4474), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
OR4X1 inst_cellmath__15__3__I11232 (.Y(N4437), .A(b_man[10]), .B(b_man[8]), .C(b_man[9]), .D(b_man[7]));
OR4X1 inst_cellmath__15__3__I11233 (.Y(N4447), .A(b_man[6]), .B(b_man[4]), .C(b_man[5]), .D(b_man[3]));
NOR2XL inst_cellmath__15__3__I861 (.Y(N4468), .A(N4464), .B(N4474));
NAND3XL inst_cellmath__15__3__I4739 (.Y(N10769), .A(N4433), .B(N4462), .C(N4468));
OR4X1 inst_cellmath__15__3__I11234 (.Y(inst_cellmath__15), .A(N4447), .B(N4437), .C(N4454), .D(N10769));
NOR2XL cynw_cm_float_add2_ieee_I865 (.Y(inst_cellmath__17), .A(inst_cellmath__14), .B(inst_cellmath__15));
XOR2XL inst_cellmath__33_49_24_I10970 (.Y(inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
NAND2BXL cynw_cm_float_add2_ieee_I4552 (.Y(inst_cellmath__13), .AN(inst_cellmath__9), .B(inst_cellmath__10));
NAND2BXL cynw_cm_float_add2_ieee_I4553 (.Y(inst_cellmath__18), .AN(inst_cellmath__14), .B(inst_cellmath__15));
NAND2XL hyperpropagate_3_1_A_I4741 (.Y(N10775), .A(inst_cellmath__18), .B(inst_cellmath__13));
AOI31X1 hyperpropagate_3_1_A_I11235 (.Y(N4525), .A0(inst_cellmath__12), .A1(inst_cellmath__39[25]), .A2(inst_cellmath__17), .B0(N10775));
INVX1 cynw_cm_float_add2_ieee_I874 (.Y(inst_cellmath__63), .A(N4525));
OR4X1 inst_cellmath__33_49_24_I11236 (.Y(N17830), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 inst_cellmath__33_49_24_I11237 (.Y(N17805), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL inst_cellmath__33_49_24_I11172 (.Y(inst_cellmath__11), .A(N17830), .B(N17805));
OR4X1 inst_cellmath__33_49_24_I11238 (.Y(N17818), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 inst_cellmath__33_49_24_I11239 (.Y(N17825), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL inst_cellmath__33_49_24_I11175 (.Y(inst_cellmath__16), .A(N17818), .B(N17825));
AND2XL cynw_cm_float_add2_ieee_I889 (.Y(N706), .A(inst_cellmath__11), .B(inst_cellmath__16));
INVXL inst_cellmath__6_0_I890 (.Y(N4581), .A(rm[0]));
INVXL inst_cellmath__6_0_I891 (.Y(N4582), .A(rm[2]));
AND3XL inst_cellmath__6_0_I4556 (.Y(inst_cellmath__6), .A(rm[1]), .B(N4582), .C(N4581));
INVX1 cynw_cm_float_add2_ieee_I15 (.Y(N556), .A(b_exp[0]));
INVX2 cynw_cm_float_add2_ieee_I16 (.Y(N557), .A(b_exp[1]));
INVX2 cynw_cm_float_add2_ieee_I17 (.Y(N558), .A(b_exp[2]));
INVX3 cynw_cm_float_add2_ieee_I18 (.Y(N559), .A(b_exp[3]));
INVX1 cynw_cm_float_add2_ieee_I19 (.Y(N560), .A(b_exp[4]));
INVX2 cynw_cm_float_add2_ieee_I20 (.Y(N561), .A(b_exp[5]));
INVX2 cynw_cm_float_add2_ieee_I21 (.Y(N562), .A(b_exp[6]));
INVX2 cynw_cm_float_add2_ieee_I22 (.Y(N563), .A(b_exp[7]));
NAND2X1 inst_cellmath__28__8__I894 (.Y(N4677), .A(a_exp[0]), .B(N556));
NOR2X1 inst_cellmath__28__8__I895 (.Y(N4594), .A(a_exp[1]), .B(N557));
NAND2X1 inst_cellmath__28__8__I896 (.Y(N4614), .A(a_exp[1]), .B(N557));
NOR2X1 inst_cellmath__28__8__I897 (.Y(N4640), .A(a_exp[2]), .B(N558));
NAND2X2 inst_cellmath__28__8__I898 (.Y(N4666), .A(a_exp[2]), .B(N558));
NOR2X1 inst_cellmath__28__8__I899 (.Y(N4687), .A(a_exp[3]), .B(N559));
NAND2X4 inst_cellmath__28__8__I900 (.Y(N4602), .A(a_exp[3]), .B(N559));
NOR2XL inst_cellmath__28__8__I901 (.Y(N4625), .A(a_exp[4]), .B(N560));
NAND2X1 inst_cellmath__28__8__I902 (.Y(N4650), .A(a_exp[4]), .B(N560));
NOR2XL inst_cellmath__28__8__I903 (.Y(N4674), .A(a_exp[5]), .B(N561));
NAND2X2 inst_cellmath__28__8__I904 (.Y(N4697), .A(a_exp[5]), .B(N561));
NOR2XL inst_cellmath__28__8__I905 (.Y(N4609), .A(a_exp[6]), .B(N562));
NAND2X1 inst_cellmath__28__8__I906 (.Y(N4635), .A(a_exp[6]), .B(N562));
NOR2XL inst_cellmath__28__8__I907 (.Y(N4659), .A(a_exp[7]), .B(N563));
NAND2X2 inst_cellmath__28__8__I908 (.Y(N4682), .A(a_exp[7]), .B(N563));
INVXL inst_cellmath__28__8__I909 (.Y(N4592), .A(N4677));
AOI21XL inst_cellmath__28__8__I910 (.Y(N4645), .A0(N4614), .A1(N4677), .B0(N4594));
INVXL inst_cellmath__28__8__I911 (.Y(N4610), .A(N4645));
AOI21XL inst_cellmath__28__8__I912 (.Y(N4692), .A0(N4666), .A1(N4594), .B0(N4640));
NAND2XL inst_cellmath__28__8__I913 (.Y(N4606), .A(N4666), .B(N4614));
AOI21X2 inst_cellmath__28__8__I914 (.Y(N4631), .A0(N4640), .A1(N4602), .B0(N4687));
NAND2X1 inst_cellmath__28__8__I915 (.Y(N4654), .A(N4602), .B(N4666));
AOI21XL inst_cellmath__28__8__I916 (.Y(N4678), .A0(N4650), .A1(N4687), .B0(N4625));
NAND2XL inst_cellmath__28__8__I917 (.Y(N4596), .A(N4650), .B(N4602));
AOI21X1 inst_cellmath__28__8__I918 (.Y(N4615), .A0(N4625), .A1(N4697), .B0(N4674));
NAND2X1 inst_cellmath__28__8__I919 (.Y(N4641), .A(N4697), .B(N4650));
AOI21XL inst_cellmath__28__8__I920 (.Y(N4668), .A0(N4635), .A1(N4674), .B0(N4609));
NAND2XL inst_cellmath__28__8__I921 (.Y(N4688), .A(N4635), .B(N4697));
AOI21X1 inst_cellmath__28__8__I922 (.Y(N4603), .A0(N4682), .A1(N4609), .B0(N4659));
NAND2X1 inst_cellmath__28__8__I923 (.Y(N4627), .A(N4682), .B(N4635));
INVXL inst_cellmath__28__8__I924 (.Y(N4662), .A(N4592));
OAI21XL inst_cellmath__28__8__I925 (.Y(N4638), .A0(N4606), .A1(N4592), .B0(N4692));
OAI21XL inst_cellmath__28__8__I927 (.Y(N4624), .A0(N4596), .A1(N4692), .B0(N4678));
NOR2XL inst_cellmath__28__8__I928 (.Y(N4648), .A(N4596), .B(N4606));
OAI21XL inst_cellmath__28__8__I929 (.Y(N4673), .A0(N4641), .A1(N4631), .B0(N4615));
NOR2XL inst_cellmath__28__8__I930 (.Y(N4695), .A(N4641), .B(N4654));
OAI21XL inst_cellmath__28__8__I931 (.Y(N4607), .A0(N4688), .A1(N4678), .B0(N4668));
NOR2XL inst_cellmath__28__8__I932 (.Y(N4634), .A(N4688), .B(N4596));
AOI21XL inst_cellmath__28__8__I935 (.Y(N4676), .A0(N4648), .A1(N4662), .B0(N4624));
AOI21XL inst_cellmath__28__8__I936 (.Y(N4613), .A0(N4695), .A1(N4610), .B0(N4673));
AOI21XL inst_cellmath__28__8__I937 (.Y(N4665), .A0(N4634), .A1(N4638), .B0(N4607));
NAND2BXL inst_cellmath__28__8__I938 (.Y(N4630), .AN(N4594), .B(N4614));
NAND2BXL inst_cellmath__28__8__I939 (.Y(N4595), .AN(N4640), .B(N4666));
NAND2BXL inst_cellmath__28__8__I940 (.Y(N4667), .AN(N4687), .B(N4602));
NAND2BXL inst_cellmath__28__8__I941 (.Y(N4626), .AN(N4625), .B(N4650));
NAND2BXL inst_cellmath__28__8__I942 (.Y(N4591), .AN(N4674), .B(N4697));
NAND2BXL inst_cellmath__28__8__I943 (.Y(N4661), .AN(N4609), .B(N4635));
NAND2BXL inst_cellmath__28__8__I944 (.Y(N4623), .AN(N4659), .B(N4682));
XNOR2X1 inst_cellmath__28__8__I945 (.Y(N565), .A(a_exp[0]), .B(N556));
XNOR2X1 inst_cellmath__28__8__I946 (.Y(N566), .A(N4662), .B(N4630));
XNOR2X1 inst_cellmath__28__8__I947 (.Y(N567), .A(N4610), .B(N4595));
OAI21XL cynw_cm_float_add2_ieee_I11038 (.Y(N4685), .A0(N4654), .A1(N4645), .B0(N4631));
XNOR2X1 inst_cellmath__28__8__I949 (.Y(N569), .A(N4685), .B(N4626));
XOR2XL inst_cellmath__28__8__I950 (.Y(N570), .A(N4676), .B(N4591));
XOR2XL inst_cellmath__28__8__I951 (.Y(N571), .A(N4613), .B(N4661));
XOR2XL inst_cellmath__28__8__I952 (.Y(N572), .A(N4665), .B(N4623));
INVXL inst_cellmath__28__8__I954 (.Y(N4643), .A(a_exp[0]));
INVXL inst_cellmath__28__8__I955 (.Y(N4690), .A(N556));
INVXL inst_cellmath__28__8__I956 (.Y(N4656), .A(N4643));
NAND2XL inst_cellmath__28__8__I957 (.Y(N4658), .A(N4690), .B(N4643));
INVXL inst_cellmath__28__8__I958 (.Y(N4619), .A(N4594));
NAND2XL inst_cellmath__28__8__I959 (.Y(N4671), .A(N4614), .B(N4690));
INVXL inst_cellmath__28__8__I961 (.Y(N4680), .A(N4656));
INVXL inst_cellmath__28__8__I962 (.Y(N4598), .A(N4658));
OAI21XL inst_cellmath__28__8__I963 (.Y(N4637), .A0(N4671), .A1(N4656), .B0(N4619));
OAI21XL inst_cellmath__28__8__I964 (.Y(N4684), .A0(N4606), .A1(N4658), .B0(N4692));
OAI21X1 inst_cellmath__28__8__I965 (.Y(N4621), .A0(N4654), .A1(N4619), .B0(N4631));
NOR2XL inst_cellmath__28__8__I966 (.Y(N4647), .A(N4654), .B(N4671));
AOI21XL inst_cellmath__28__8__I969 (.Y(N4611), .A0(N4647), .A1(N4680), .B0(N4621));
AOI21XL inst_cellmath__28__8__I970 (.Y(N4664), .A0(N4648), .A1(N4598), .B0(N4624));
AOI21XL inst_cellmath__28__8__I971 (.Y(N4601), .A0(N4695), .A1(N4637), .B0(N4673));
AOI21XL inst_cellmath__28__8__I972 (.Y(N4649), .A0(N4634), .A1(N4684), .B0(N4607));
INVXL cynw_cm_float_add2_ieee_I11042 (.Y(N4617), .A(N4680));
XOR2XL inst_cellmath__28__8__I976 (.Y(inst_cellmath__27[0]), .A(N4617), .B(N4690));
XOR2XL inst_cellmath__28__8__I977 (.Y(inst_cellmath__27[1]), .A(N4598), .B(N4630));
XOR2XL inst_cellmath__28__8__I978 (.Y(inst_cellmath__27[2]), .A(N4637), .B(N4595));
XNOR2X1 inst_cellmath__28__8__I980 (.Y(inst_cellmath__27[4]), .A(N4611), .B(N4626));
XNOR2X1 inst_cellmath__28__8__I981 (.Y(inst_cellmath__27[5]), .A(N4664), .B(N4591));
XNOR2X1 inst_cellmath__28__8__I982 (.Y(inst_cellmath__27[6]), .A(N4601), .B(N4661));
CLKINVX8 inst_cellmath__34_0_I985 (.Y(N4820), .A(a_man[1]));
CLKINVX6 inst_cellmath__34_0_I987 (.Y(N4801), .A(a_man[3]));
INVX3 inst_cellmath__34_0_I988 (.Y(N4866), .A(a_man[4]));
CLKINVX4 inst_cellmath__34_0_I989 (.Y(N4934), .A(a_man[5]));
CLKINVX4 inst_cellmath__34_0_I990 (.Y(N4847), .A(a_man[6]));
CLKINVX8 inst_cellmath__34_0_I991 (.Y(N4912), .A(a_man[7]));
INVX2 inst_cellmath__34_0_I992 (.Y(N4829), .A(a_man[8]));
INVX3 inst_cellmath__34_0_I993 (.Y(N4893), .A(a_man[9]));
INVX1 inst_cellmath__34_0_I994 (.Y(N4807), .A(a_man[10]));
CLKINVX4 inst_cellmath__34_0_I995 (.Y(N4875), .A(a_man[11]));
INVX2 inst_cellmath__34_0_I996 (.Y(N4791), .A(a_man[12]));
CLKINVX6 inst_cellmath__34_0_I997 (.Y(N4854), .A(a_man[13]));
INVX2 inst_cellmath__34_0_I998 (.Y(N4922), .A(a_man[14]));
CLKINVX6 inst_cellmath__34_0_I999 (.Y(N4839), .A(a_man[15]));
INVX1 inst_cellmath__34_0_I1000 (.Y(N4901), .A(a_man[16]));
INVX2 inst_cellmath__34_0_I1001 (.Y(N4817), .A(a_man[17]));
INVXL inst_cellmath__34_0_I1002 (.Y(N4884), .A(a_man[18]));
INVX2 inst_cellmath__34_0_I1003 (.Y(N4796), .A(a_man[19]));
INVX2 inst_cellmath__34_0_I1004 (.Y(N4864), .A(a_man[20]));
INVX2 inst_cellmath__34_0_I1005 (.Y(N4931), .A(a_man[21]));
INVX1 inst_cellmath__34_0_I1006 (.Y(N4843), .A(a_man[22]));
NAND2X4 inst_cellmath__34_0_I1007 (.Y(N4835), .A(b_man[1]), .B(N4820));
NOR2X4 inst_cellmath__34_0_I1008 (.Y(N4800), .A(b_man[1]), .B(N4820));
NAND2X1 inst_cellmath__34_0_I1009 (.Y(N4933), .A(b_man[2]), .B(N4338));
NOR2X1 inst_cellmath__34_0_I1010 (.Y(N4898), .A(b_man[2]), .B(N4338));
NAND2X1 inst_cellmath__34_0_I1011 (.Y(N4880), .A(b_man[3]), .B(N4801));
NOR2X4 inst_cellmath__34_0_I1012 (.Y(N4846), .A(b_man[3]), .B(N4801));
NAND2X2 inst_cellmath__34_0_I1013 (.Y(N4828), .A(b_man[4]), .B(N4866));
NOR2XL inst_cellmath__34_0_I1014 (.Y(N4794), .A(b_man[4]), .B(N4866));
NAND2X1 inst_cellmath__34_0_I1015 (.Y(N4927), .A(b_man[5]), .B(N4934));
NOR2X4 inst_cellmath__34_0_I1016 (.Y(N4892), .A(b_man[5]), .B(N4934));
NAND2XL inst_cellmath__34_0_I1017 (.Y(N4874), .A(b_man[6]), .B(N4847));
NOR2X2 inst_cellmath__34_0_I1018 (.Y(N4841), .A(b_man[6]), .B(N4847));
NAND2X1 inst_cellmath__34_0_I1019 (.Y(N4823), .A(b_man[7]), .B(N4912));
NOR2X6 inst_cellmath__34_0_I1020 (.Y(N4790), .A(b_man[7]), .B(N4912));
NAND2X2 inst_cellmath__34_0_I1021 (.Y(N4921), .A(b_man[8]), .B(N4829));
NOR2XL inst_cellmath__34_0_I1022 (.Y(N4889), .A(b_man[8]), .B(N4829));
NAND2X1 inst_cellmath__34_0_I1023 (.Y(N4869), .A(b_man[9]), .B(N4893));
NOR2X4 inst_cellmath__34_0_I1024 (.Y(N4837), .A(b_man[9]), .B(N4893));
NAND2XL inst_cellmath__34_0_I1025 (.Y(N4816), .A(b_man[10]), .B(N4807));
NAND2XL inst_cellmath__34_0_I1027 (.Y(N4915), .A(b_man[11]), .B(N4875));
NOR2X4 inst_cellmath__34_0_I1028 (.Y(N4882), .A(b_man[11]), .B(N4875));
NAND2XL inst_cellmath__34_0_I1029 (.Y(N4863), .A(b_man[12]), .B(N4791));
NOR2XL inst_cellmath__34_0_I1030 (.Y(N4832), .A(b_man[12]), .B(N4791));
NAND2X1 inst_cellmath__34_0_I1031 (.Y(N4810), .A(b_man[13]), .B(N4854));
NOR2X6 inst_cellmath__34_0_I1032 (.Y(N4929), .A(b_man[13]), .B(N4854));
NAND2XL inst_cellmath__34_0_I1033 (.Y(N4910), .A(b_man[14]), .B(N4922));
NOR2X2 inst_cellmath__34_0_I1034 (.Y(N4878), .A(b_man[14]), .B(N4922));
NAND2X1 inst_cellmath__34_0_I1035 (.Y(N4857), .A(b_man[15]), .B(N4839));
NOR2X4 inst_cellmath__34_0_I1036 (.Y(N4825), .A(b_man[15]), .B(N4839));
NAND2XL inst_cellmath__34_0_I1037 (.Y(N4805), .A(b_man[16]), .B(N4901));
NOR2XL inst_cellmath__34_0_I1038 (.Y(N4924), .A(b_man[16]), .B(N4901));
NAND2XL inst_cellmath__34_0_I1039 (.Y(N4904), .A(b_man[17]), .B(N4817));
NOR2X2 inst_cellmath__34_0_I1040 (.Y(N4871), .A(b_man[17]), .B(N4817));
NAND2XL inst_cellmath__34_0_I1041 (.Y(N4851), .A(b_man[18]), .B(N4884));
NOR2XL inst_cellmath__34_0_I1042 (.Y(N4819), .A(b_man[18]), .B(N4884));
NAND2XL inst_cellmath__34_0_I1043 (.Y(N4799), .A(b_man[19]), .B(N4796));
NOR2X2 inst_cellmath__34_0_I1044 (.Y(N4917), .A(b_man[19]), .B(N4796));
NAND2XL inst_cellmath__34_0_I1045 (.Y(N4897), .A(b_man[20]), .B(N4864));
NOR2X1 inst_cellmath__34_0_I1046 (.Y(N4865), .A(b_man[20]), .B(N4864));
NAND2XL inst_cellmath__34_0_I1047 (.Y(N4845), .A(b_man[21]), .B(N4931));
NOR2X1 inst_cellmath__34_0_I1048 (.Y(N4812), .A(b_man[21]), .B(N4931));
AND2XL inst_cellmath__34_0_I1049 (.Y(N4830), .A(b_man[22]), .B(N4843));
OR2XL inst_cellmath__34_0_I1050 (.Y(N4861), .A(b_man[22]), .B(N4843));
OAI21XL inst_cellmath__34_0_I1051 (.Y(N4859), .A0(N4897), .A1(N4812), .B0(N4845));
NOR2X1 inst_cellmath__34_0_I1052 (.Y(N4891), .A(N4865), .B(N4812));
OAI21X1 inst_cellmath__34_0_I1053 (.Y(N4926), .A0(N4917), .A1(N4851), .B0(N4799));
NOR2X1 inst_cellmath__34_0_I1054 (.Y(N4806), .A(N4917), .B(N4819));
OAI21X1 inst_cellmath__34_0_I1055 (.Y(N4840), .A0(N4871), .A1(N4805), .B0(N4904));
NOR2XL inst_cellmath__34_0_I1056 (.Y(N4873), .A(N4871), .B(N4924));
OAI21X2 inst_cellmath__34_0_I1057 (.Y(N4906), .A0(N4825), .A1(N4910), .B0(N4857));
NOR2X2 inst_cellmath__34_0_I1058 (.Y(N4789), .A(N4878), .B(N4825));
OAI21X2 inst_cellmath__34_0_I1059 (.Y(N4822), .A0(N4929), .A1(N4863), .B0(N4810));
NOR2X1 inst_cellmath__34_0_I1060 (.Y(N4853), .A(N4832), .B(N4929));
OAI21X1 inst_cellmath__34_0_I1061 (.Y(N4888), .A0(N4882), .A1(N4816), .B0(N4915));
AOI2BB1X1 inst_cellmath__34_0_I4558 (.Y(N4919), .A0N(b_man[10]), .A1N(N4807), .B0(N4882));
OAI21X2 inst_cellmath__34_0_I1063 (.Y(N4802), .A0(N4921), .A1(N4837), .B0(N4869));
NOR2XL inst_cellmath__34_0_I1064 (.Y(N4836), .A(N4889), .B(N4837));
OAI21X2 inst_cellmath__34_0_I1065 (.Y(N4868), .A0(N4790), .A1(N4874), .B0(N4823));
NOR2X1 inst_cellmath__34_0_I1066 (.Y(N4899), .A(N4841), .B(N4790));
OAI21X2 inst_cellmath__34_0_I1067 (.Y(N4935), .A0(N4828), .A1(N4892), .B0(N4927));
NOR2XL inst_cellmath__34_0_I1068 (.Y(N4814), .A(N4892), .B(N4794));
OAI21X2 inst_cellmath__34_0_I1069 (.Y(N4848), .A0(N4846), .A1(N4933), .B0(N4880));
NOR2XL inst_cellmath__34_0_I1070 (.Y(N4881), .A(N4898), .B(N4846));
CLKINVX4 inst_cellmath__34_0_I1071 (.Y(N4911), .A(b_man[0]));
OAI31X4 inst_cellmath__34_0_I1072 (.Y(N4914), .A0(N4911), .A1(a_man[0]), .A2(N4800), .B0(N4835));
AOI21XL inst_cellmath__34_0_I1073 (.Y(N4894), .A0(N4861), .A1(N4859), .B0(N4830));
NAND2X1 inst_cellmath__34_0_I1074 (.Y(N4928), .A(N4861), .B(N4891));
AOI21X1 inst_cellmath__34_0_I1075 (.Y(N4809), .A0(N4806), .A1(N4840), .B0(N4926));
AOI21X2 inst_cellmath__34_0_I1076 (.Y(N4876), .A0(N4789), .A1(N4822), .B0(N4906));
NAND2X1 inst_cellmath__34_0_I1077 (.Y(N4908), .A(N4789), .B(N4853));
AOI21X1 inst_cellmath__34_0_I1078 (.Y(N4792), .A0(N4802), .A1(N4919), .B0(N4888));
NAND2XL inst_cellmath__34_0_I1079 (.Y(N4824), .A(N4836), .B(N4919));
AOI21X1 inst_cellmath__34_0_I1080 (.Y(N4856), .A0(N4899), .A1(N4935), .B0(N4868));
NAND2XL inst_cellmath__34_0_I1081 (.Y(N4890), .A(N4899), .B(N4814));
AOI21X1 inst_cellmath__34_0_I1082 (.Y(N4923), .A0(N4881), .A1(N4914), .B0(N4848));
OAI21X1 inst_cellmath__34_0_I1084 (.Y(N4903), .A0(N4908), .A1(N4792), .B0(N4876));
NOR2XL inst_cellmath__34_0_I1085 (.Y(N4938), .A(N4908), .B(N4824));
OAI21X2 inst_cellmath__34_0_I1086 (.Y(N4818), .A0(N4890), .A1(N4923), .B0(N4856));
OAI21X1 cynw_cm_float_add2_ieee_I11039 (.Y(N17588), .A0(N4627), .A1(N4615), .B0(N4603));
NOR2X1 cynw_cm_float_add2_ieee_I11040 (.Y(N17597), .A(N4627), .B(N4641));
AO21X1 cynw_cm_float_add2_ieee_I11041 (.Y(N573), .A0(N17597), .A1(N4685), .B0(N17588));
AOI21X2 cynw_cm_float_add2_ieee_I11043 (.Y(N17583), .A0(N17597), .A1(N4621), .B0(N17588));
NAND2X2 cynw_cm_float_add2_ieee_I11044 (.Y(N17592), .A(N17597), .B(N4647));
NOR2X1 cynw_cm_float_add2_ieee_I11045 (.Y(N17569), .A(N4617), .B(N17592));
INVX1 cynw_cm_float_add2_ieee_I11046 (.Y(N17576), .A(N17583));
NOR2X4 cynw_cm_float_add2_ieee_I11047 (.Y(N17590), .A(N17569), .B(N17576));
XOR2XL cynw_cm_float_add2_ieee_I11186 (.Y(N17859), .A(N4638), .B(N4667));
XNOR2X1 cynw_cm_float_add2_ieee_I11187 (.Y(N17869), .A(N4684), .B(N4667));
OAI21X4 cynw_cm_float_add2_ieee_I11188 (.Y(inst_cellmath__27[8]), .A0(N17592), .A1(N4617), .B0(N17583));
MX2XL cynw_cm_float_add2_ieee_I11189 (.Y(inst_cellmath__35[1]), .A(inst_cellmath__27[1]), .B(N566), .S0(inst_cellmath__27[8]));
MXI2XL cynw_cm_float_add2_ieee_I11253 (.Y(inst_cellmath__35[3]), .A(N17869), .B(N17859), .S0(inst_cellmath__27[8]));
INVXL cynw_cm_float_add2_ieee_I1155 (.Y(N5206), .A(b_man[13]));
NAND3BX1 cynw_cm_float_add2_ieee_I11049 (.Y(N17571), .AN(N4928), .B(N4806), .C(N4873));
AOI21X2 cynw_cm_float_add2_ieee_I11050 (.Y(N17578), .A0(N4938), .A1(N4818), .B0(N4903));
OA21X1 cynw_cm_float_add2_ieee_I11051 (.Y(N17586), .A0(N4928), .A1(N4809), .B0(N4894));
OAI21X4 cynw_cm_float_add2_ieee_I11052 (.Y(N17595), .A0(N17571), .A1(N17578), .B0(N17586));
NAND2X4 cynw_cm_float_add2_ieee_I11053 (.Y(N17580), .A(N573), .B(N17595));
NAND2X8 cynw_cm_float_add2_ieee_I11054 (.Y(N4309), .A(N17590), .B(N17580));
MXI2XL cynw_cm_float_add2_ieee_I1184 (.Y(inst_cellmath__36[39]), .A(N5206), .B(N4854), .S0(N4309));
INVXL cynw_cm_float_add2_ieee_I1154 (.Y(N5180), .A(b_man[12]));
MXI2XL cynw_cm_float_add2_ieee_I1183 (.Y(inst_cellmath__36[38]), .A(N5180), .B(N4791), .S0(N4309));
MXI2X4 inst_cellmath__37_0_I4326 (.Y(N5376), .A(inst_cellmath__27[0]), .B(N565), .S0(inst_cellmath__27[8]));
MX2XL cynw_cm_float_add2_ieee_I11192 (.Y(N5412), .A(inst_cellmath__36[39]), .B(inst_cellmath__36[38]), .S0(N5376));
INVXL cynw_cm_float_add2_ieee_I1157 (.Y(N5259), .A(b_man[15]));
MXI2XL cynw_cm_float_add2_ieee_I1186 (.Y(inst_cellmath__36[41]), .A(N5259), .B(N4839), .S0(N4309));
INVXL cynw_cm_float_add2_ieee_I1156 (.Y(N5233), .A(b_man[14]));
MXI2XL cynw_cm_float_add2_ieee_I1185 (.Y(inst_cellmath__36[40]), .A(N5233), .B(N4922), .S0(N4309));
MX2XL cynw_cm_float_add2_ieee_I11193 (.Y(N5519), .A(inst_cellmath__36[41]), .B(inst_cellmath__36[40]), .S0(N5376));
INVXL cynw_cm_float_add2_ieee_I1159 (.Y(N5191), .A(b_man[17]));
MXI2XL cynw_cm_float_add2_ieee_I1188 (.Y(inst_cellmath__36[43]), .A(N5191), .B(N4817), .S0(N4309));
INVXL cynw_cm_float_add2_ieee_I1158 (.Y(N5164), .A(b_man[16]));
MXI2XL cynw_cm_float_add2_ieee_I1187 (.Y(inst_cellmath__36[42]), .A(N5164), .B(N4901), .S0(N4309));
MX2XL cynw_cm_float_add2_ieee_I11194 (.Y(N5379), .A(inst_cellmath__36[43]), .B(inst_cellmath__36[42]), .S0(N5376));
INVXL cynw_cm_float_add2_ieee_I1161 (.Y(N5244), .A(b_man[19]));
MXI2XL cynw_cm_float_add2_ieee_I1190 (.Y(inst_cellmath__36[45]), .A(N5244), .B(N4796), .S0(N4309));
INVXL cynw_cm_float_add2_ieee_I1160 (.Y(N5217), .A(b_man[18]));
MXI2XL cynw_cm_float_add2_ieee_I1189 (.Y(inst_cellmath__36[44]), .A(N5217), .B(N4884), .S0(N4309));
MX2XL cynw_cm_float_add2_ieee_I11195 (.Y(N5486), .A(inst_cellmath__36[45]), .B(inst_cellmath__36[44]), .S0(N5376));
INVXL cynw_cm_float_add2_ieee_I1163 (.Y(N5175), .A(b_man[21]));
MXI2XL cynw_cm_float_add2_ieee_I1192 (.Y(inst_cellmath__36[47]), .A(N5175), .B(N4931), .S0(N4309));
INVXL cynw_cm_float_add2_ieee_I1162 (.Y(N5148), .A(b_man[20]));
MXI2XL cynw_cm_float_add2_ieee_I1191 (.Y(inst_cellmath__36[46]), .A(N5148), .B(N4864), .S0(N4309));
MX2XL cynw_cm_float_add2_ieee_I11196 (.Y(N5346), .A(inst_cellmath__36[47]), .B(inst_cellmath__36[46]), .S0(N5376));
INVXL cynw_cm_float_add2_ieee_I1164 (.Y(N5201), .A(b_man[22]));
MXI2XL cynw_cm_float_add2_ieee_I1193 (.Y(inst_cellmath__36[48]), .A(N5201), .B(N4843), .S0(N4309));
NAND2BXL cynw_cm_float_add2_ieee_I11197 (.Y(N5454), .AN(inst_cellmath__36[48]), .B(N5376));
MX2XL inst_cellmath__35_0_I1106 (.Y(inst_cellmath__35[2]), .A(inst_cellmath__27[2]), .B(N567), .S0(inst_cellmath__27[8]));
CLKINVX12 cynw_cm_float_add2_ieee_I11198 (.Y(N5560), .A(inst_cellmath__35[2]));
MXI2X1 cynw_cm_float_add2_ieee_I11199 (.Y(N5461), .A(N5379), .B(N5412), .S0(N5560));
INVX1 cynw_cm_float_add2_ieee_I11200 (.Y(N17895), .A(N5560));
MXI2X1 cynw_cm_float_add2_ieee_I11201 (.Y(N5571), .A(N5519), .B(N5486), .S0(N17895));
INVXL cynw_cm_float_add2_ieee_I11202 (.Y(N17851), .A(N17895));
NAND2XL cynw_cm_float_add2_ieee_I11203 (.Y(N5398), .A(N17851), .B(N5346));
NAND2XL cynw_cm_float_add2_ieee_I11204 (.Y(N5367), .A(N17851), .B(N5454));
BUFX6 cynw_cm_float_add2_ieee_I11205 (.Y(N5496), .A(inst_cellmath__35[1]));
MXI2X1 cynw_cm_float_add2_ieee_I11206 (.Y(N5459), .A(N5461), .B(N5571), .S0(N5496));
MXI2XL cynw_cm_float_add2_ieee_I11207 (.Y(N5396), .A(N5398), .B(N5367), .S0(N5496));
INVX2 cynw_cm_float_add2_ieee_I11208 (.Y(N5347), .A(inst_cellmath__35[3]));
MXI2XL cynw_cm_float_add2_ieee_I11209 (.Y(N5426), .A(N5396), .B(N5459), .S0(N5347));
MX2XL cynw_cm_float_add2_ieee_I1095 (.Y(inst_cellmath__48), .A(a_sign), .B(b_sign), .S0(N4309));
XNOR2X1 inst_cellmath__35_0_I4345 (.Y(N5094), .A(N4649), .B(N4623));
MX2XL inst_cellmath__35_0_I1108 (.Y(inst_cellmath__35[4]), .A(inst_cellmath__27[4]), .B(N569), .S0(inst_cellmath__27[8]));
MX2XL inst_cellmath__35_0_I1109 (.Y(inst_cellmath__35[5]), .A(inst_cellmath__27[5]), .B(N570), .S0(inst_cellmath__27[8]));
MX2XL inst_cellmath__35_0_I1110 (.Y(inst_cellmath__35[6]), .A(inst_cellmath__27[6]), .B(N571), .S0(inst_cellmath__27[8]));
MX2XL inst_cellmath__35_0_I1111 (.Y(inst_cellmath__35[7]), .A(N5094), .B(N572), .S0(inst_cellmath__27[8]));
NOR2XL inst_cellmath__30_0_I1112 (.Y(N5114), .A(inst_cellmath__35[2]), .B(inst_cellmath__35[1]));
NAND2XL inst_cellmath__30_0_I1113 (.Y(N5119), .A(inst_cellmath__35[3]), .B(inst_cellmath__35[4]));
NOR3XL inst_cellmath__30_0_I1114 (.Y(N5123), .A(inst_cellmath__35[7]), .B(inst_cellmath__35[6]), .C(inst_cellmath__35[5]));
OAI21X1 inst_cellmath__30_0_I1115 (.Y(inst_cellmath__30), .A0(N5114), .A1(N5119), .B0(N5123));
INVXL cynw_cm_float_add2_ieee_I1119 (.Y(N5224), .A(a_man[0]));
INVXL cynw_cm_float_add2_ieee_I1143 (.Y(N5253), .A(b_man[1]));
INVXL cynw_cm_float_add2_ieee_I1145 (.Y(N5184), .A(b_man[3]));
INVXL cynw_cm_float_add2_ieee_I1146 (.Y(N5210), .A(b_man[4]));
INVXL cynw_cm_float_add2_ieee_I1147 (.Y(N5237), .A(b_man[5]));
INVXL cynw_cm_float_add2_ieee_I1148 (.Y(N5141), .A(b_man[6]));
INVXL cynw_cm_float_add2_ieee_I1149 (.Y(N5168), .A(b_man[7]));
INVXL cynw_cm_float_add2_ieee_I1150 (.Y(N5195), .A(b_man[8]));
INVXL cynw_cm_float_add2_ieee_I1151 (.Y(N5222), .A(b_man[9]));
INVXL cynw_cm_float_add2_ieee_I1152 (.Y(N5249), .A(b_man[10]));
INVXL cynw_cm_float_add2_ieee_I1153 (.Y(N5153), .A(b_man[11]));
MXI2XL cynw_cm_float_add2_ieee_I1171 (.Y(inst_cellmath__36[26]), .A(N4911), .B(N5224), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1172 (.Y(inst_cellmath__36[27]), .A(N5253), .B(N4820), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1173 (.Y(inst_cellmath__36[28]), .A(N4433), .B(N4338), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1174 (.Y(inst_cellmath__36[29]), .A(N5184), .B(N4801), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1175 (.Y(inst_cellmath__36[30]), .A(N5210), .B(N4866), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1176 (.Y(inst_cellmath__36[31]), .A(N5237), .B(N4934), .S0(N4309));
MXI2X1 cynw_cm_float_add2_ieee_I1177 (.Y(inst_cellmath__36[32]), .A(N5141), .B(N4847), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1178 (.Y(inst_cellmath__36[33]), .A(N5168), .B(N4912), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1179 (.Y(inst_cellmath__36[34]), .A(N5195), .B(N4829), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1180 (.Y(inst_cellmath__36[35]), .A(N5222), .B(N4893), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1181 (.Y(inst_cellmath__36[36]), .A(N5249), .B(N4807), .S0(N4309));
MXI2XL cynw_cm_float_add2_ieee_I1182 (.Y(inst_cellmath__36[37]), .A(N5153), .B(N4875), .S0(N4309));
NOR2BX1 inst_cellmath__37_0_I1202 (.Y(N5397), .AN(inst_cellmath__36[26]), .B(N5376));
MX2XL inst_cellmath__37_0_I1203 (.Y(N5505), .A(inst_cellmath__36[27]), .B(inst_cellmath__36[26]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1204 (.Y(N5559), .A(inst_cellmath__36[28]), .B(inst_cellmath__36[27]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1205 (.Y(N5366), .A(inst_cellmath__36[29]), .B(inst_cellmath__36[28]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1206 (.Y(N5420), .A(inst_cellmath__36[30]), .B(inst_cellmath__36[29]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1207 (.Y(N5473), .A(inst_cellmath__36[31]), .B(inst_cellmath__36[30]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1208 (.Y(N5527), .A(inst_cellmath__36[32]), .B(inst_cellmath__36[31]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1209 (.Y(N5583), .A(inst_cellmath__36[33]), .B(inst_cellmath__36[32]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1210 (.Y(N5387), .A(inst_cellmath__36[34]), .B(inst_cellmath__36[33]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1211 (.Y(N5443), .A(inst_cellmath__36[35]), .B(inst_cellmath__36[34]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1212 (.Y(N5495), .A(inst_cellmath__36[36]), .B(inst_cellmath__36[35]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1213 (.Y(N5551), .A(inst_cellmath__36[37]), .B(inst_cellmath__36[36]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1214 (.Y(N5355), .A(inst_cellmath__36[38]), .B(inst_cellmath__36[37]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1216 (.Y(N5464), .A(inst_cellmath__36[40]), .B(inst_cellmath__36[39]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1218 (.Y(N5574), .A(inst_cellmath__36[42]), .B(inst_cellmath__36[41]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1220 (.Y(N5434), .A(inst_cellmath__36[44]), .B(inst_cellmath__36[43]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1222 (.Y(N5541), .A(inst_cellmath__36[46]), .B(inst_cellmath__36[45]), .S0(N5376));
MX2XL inst_cellmath__37_0_I1224 (.Y(N5401), .A(inst_cellmath__36[48]), .B(inst_cellmath__36[47]), .S0(N5376));
NAND2BXL inst_cellmath__37_0_I1234 (.Y(N5568), .AN(N5560), .B(N5397));
NAND2BXL inst_cellmath__37_0_I1235 (.Y(N5428), .AN(N5560), .B(N5505));
NAND2BXL inst_cellmath__37_0_I1236 (.Y(N5535), .AN(N5560), .B(N5559));
NAND2BXL inst_cellmath__37_0_I1237 (.Y(N5395), .AN(N5560), .B(N5366));
MXI2XL inst_cellmath__37_0_I1238 (.Y(N5503), .A(N5420), .B(N5397), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1239 (.Y(N5558), .A(N5473), .B(N5505), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1240 (.Y(N5363), .A(N5527), .B(N5559), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1241 (.Y(N5418), .A(N5583), .B(N5366), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1242 (.Y(N5471), .A(N5387), .B(N5420), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1243 (.Y(N5525), .A(N5443), .B(N5473), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1244 (.Y(N5581), .A(N5495), .B(N5527), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1245 (.Y(N5385), .A(N5551), .B(N5583), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1246 (.Y(N5441), .A(N5355), .B(N5387), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1247 (.Y(N5492), .A(N5412), .B(N5443), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1248 (.Y(N5548), .A(N5464), .B(N5495), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1249 (.Y(N5352), .A(N5519), .B(N5551), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1250 (.Y(N5409), .A(N5574), .B(N5355), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1252 (.Y(N5515), .A(N5434), .B(N5464), .S0(N5560));
MXI2X1 inst_cellmath__37_0_I1254 (.Y(N5375), .A(N5541), .B(N5574), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1255 (.Y(N5431), .A(N5346), .B(N5379), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1256 (.Y(N5482), .A(N5401), .B(N5434), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1257 (.Y(N5538), .A(N5454), .B(N5486), .S0(N5560));
MXI2XL inst_cellmath__37_0_I1258 (.Y(N5342), .A(N5376), .B(N5541), .S0(N5560));
NAND2XL inst_cellmath__37_0_I1260 (.Y(N5506), .A(N5401), .B(N5560));
NAND2XL inst_cellmath__37_0_I1262 (.Y(N5474), .A(N5376), .B(N5560));
NOR2BX1 inst_cellmath__37_0_I1271 (.Y(N5563), .AN(N5496), .B(N5568));
NOR2BX1 inst_cellmath__37_0_I1272 (.Y(N5424), .AN(N5496), .B(N5428));
MXI2XL inst_cellmath__37_0_I1273 (.Y(N5531), .A(N5568), .B(N5535), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1274 (.Y(N5336), .A(N5428), .B(N5395), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1275 (.Y(N5391), .A(N5535), .B(N5503), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1276 (.Y(N5447), .A(N5395), .B(N5558), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1277 (.Y(N5499), .A(N5503), .B(N5363), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1278 (.Y(N5555), .A(N5558), .B(N5418), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1279 (.Y(N5359), .A(N5363), .B(N5471), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1280 (.Y(N5416), .A(N5418), .B(N5525), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1281 (.Y(N5468), .A(N5471), .B(N5581), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1282 (.Y(N5523), .A(N5525), .B(N5385), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1283 (.Y(N5578), .A(N5581), .B(N5441), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1284 (.Y(N5383), .A(N5385), .B(N5492), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1285 (.Y(N5438), .A(N5441), .B(N5548), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1286 (.Y(N5490), .A(N5492), .B(N5352), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1287 (.Y(N5545), .A(N5548), .B(N5409), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1288 (.Y(N5350), .A(N5352), .B(N5461), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1289 (.Y(N5406), .A(N5409), .B(N5515), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1291 (.Y(N5513), .A(N5515), .B(N5375), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1292 (.Y(N5569), .A(N5571), .B(N5431), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1293 (.Y(N5373), .A(N5375), .B(N5482), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1294 (.Y(N5429), .A(N5431), .B(N5538), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1295 (.Y(N5480), .A(N5482), .B(N5342), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1296 (.Y(N5536), .A(N5538), .B(N5398), .S0(N5496));
MXI2X1 inst_cellmath__37_0_I1297 (.Y(N5340), .A(N5342), .B(N5506), .S0(N5496));
MXI2XL inst_cellmath__37_0_I1299 (.Y(N5450), .A(N5506), .B(N5474), .S0(N5496));
NOR2XL inst_cellmath__37_0_I1300 (.Y(N5504), .A(N5367), .B(N5496));
NOR2XL inst_cellmath__37_0_I1301 (.Y(N5365), .A(N5474), .B(N5496));
NAND2BXL inst_cellmath__37_0_I1313 (.Y(N5518), .AN(N5347), .B(N5563));
NAND2BXL inst_cellmath__37_0_I1314 (.Y(N5377), .AN(N5347), .B(N5424));
NAND2BXL inst_cellmath__37_0_I1315 (.Y(N5485), .AN(N5347), .B(N5531));
NAND2BXL inst_cellmath__37_0_I1316 (.Y(N5345), .AN(N5347), .B(N5336));
NAND2BXL inst_cellmath__37_0_I1317 (.Y(N5452), .AN(N5347), .B(N5391));
NAND2BX1 inst_cellmath__37_0_I1318 (.Y(N5562), .AN(N5347), .B(N5447));
NAND2BXL inst_cellmath__37_0_I1319 (.Y(N5423), .AN(N5347), .B(N5499));
NAND2BXL inst_cellmath__37_0_I1320 (.Y(N5529), .AN(N5347), .B(N5555));
MXI2XL inst_cellmath__37_0_I1321 (.Y(N5390), .A(N5359), .B(N5563), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1322 (.Y(N5445), .A(N5416), .B(N5424), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1323 (.Y(N5498), .A(N5468), .B(N5531), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1324 (.Y(N5554), .A(N5523), .B(N5336), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1325 (.Y(N5357), .A(N5578), .B(N5391), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1326 (.Y(N5415), .A(N5383), .B(N5447), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1327 (.Y(N5467), .A(N5438), .B(N5499), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1328 (.Y(N5521), .A(N5490), .B(N5555), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1329 (.Y(N5577), .A(N5545), .B(N5359), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1330 (.Y(N5382), .A(N5350), .B(N5416), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1331 (.Y(N5436), .A(N5406), .B(N5468), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1332 (.Y(N5489), .A(N5459), .B(N5523), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1333 (.Y(N5544), .A(N5513), .B(N5578), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1334 (.Y(N5348), .A(N5569), .B(N5383), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1335 (.Y(N5405), .A(N5373), .B(N5438), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1336 (.Y(N5458), .A(N5429), .B(N5490), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1337 (.Y(N5511), .A(N5480), .B(N5545), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1338 (.Y(N5567), .A(N5536), .B(N5350), .S0(N5347));
MXI2X1 inst_cellmath__37_0_I1339 (.Y(N5372), .A(N5340), .B(N5406), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1341 (.Y(N5479), .A(N5450), .B(N5513), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1342 (.Y(N5534), .A(N5504), .B(N5569), .S0(N5347));
MXI2XL inst_cellmath__37_0_I1343 (.Y(N5338), .A(N5365), .B(N5373), .S0(N5347));
NAND2XL inst_cellmath__37_0_I1344 (.Y(N5394), .A(N5429), .B(N5347));
NAND2XL inst_cellmath__37_0_I1345 (.Y(N5501), .A(N5347), .B(N5480));
NAND2XL inst_cellmath__37_0_I1346 (.Y(N5362), .A(N5536), .B(N5347));
NAND2XL inst_cellmath__37_0_I1347 (.Y(N5470), .A(N5340), .B(N5347));
NAND2XL inst_cellmath__37_0_I1348 (.Y(N5579), .A(N5396), .B(N5347));
NAND2X1 inst_cellmath__37_0_I1349 (.Y(N5440), .A(N5347), .B(N5450));
NAND2XL inst_cellmath__37_0_I1350 (.Y(N5547), .A(N5504), .B(N5347));
NAND2X1 inst_cellmath__37_0_I1351 (.Y(N5407), .A(N5347), .B(N5365));
BUFX16 inst_cellmath__37_0_I4564 (.Y(N5360), .A(inst_cellmath__35[4]));
NOR2BX1 inst_cellmath__37_0_I1366 (.Y(inst_cellmath__37[0]), .AN(N5360), .B(N5562));
NOR2BX1 inst_cellmath__37_0_I1367 (.Y(inst_cellmath__37[1]), .AN(N5360), .B(N5423));
NOR2BX1 inst_cellmath__37_0_I1368 (.Y(inst_cellmath__37[2]), .AN(N5360), .B(N5529));
NOR2BXL inst_cellmath__37_0_I1369 (.Y(inst_cellmath__37[3]), .AN(N5360), .B(N5390));
NOR2BXL inst_cellmath__37_0_I1370 (.Y(inst_cellmath__37[4]), .AN(N5360), .B(N5445));
NOR2BXL inst_cellmath__37_0_I1371 (.Y(inst_cellmath__37[5]), .AN(N5360), .B(N5498));
NOR2BXL inst_cellmath__37_0_I1372 (.Y(inst_cellmath__37[6]), .AN(N5360), .B(N5554));
NOR2BX1 inst_cellmath__37_0_I1373 (.Y(inst_cellmath__37[7]), .AN(N5360), .B(N5357));
NOR2BX1 inst_cellmath__37_0_I1374 (.Y(inst_cellmath__37[8]), .AN(N5360), .B(N5415));
NOR2BX1 inst_cellmath__37_0_I1375 (.Y(inst_cellmath__37[9]), .AN(N5360), .B(N5467));
NOR2BXL inst_cellmath__37_0_I1376 (.Y(inst_cellmath__37[10]), .AN(N5360), .B(N5521));
MXI2XL inst_cellmath__37_0_I1377 (.Y(inst_cellmath__37[11]), .A(N5518), .B(N5577), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1378 (.Y(inst_cellmath__37[12]), .A(N5377), .B(N5382), .S0(N5360));
MXI2X1 inst_cellmath__37_0_I1379 (.Y(inst_cellmath__37[13]), .A(N5485), .B(N5436), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1380 (.Y(inst_cellmath__37[14]), .A(N5345), .B(N5489), .S0(N5360));
INVXL mx2i_A_I11452 (.Y(N17945), .A(N5360));
AOI22XL mx2i_A_I11453 (.Y(inst_cellmath__37[15]), .A0(N17945), .A1(N5452), .B0(N5544), .B1(N5360));
MXI2X1 inst_cellmath__37_0_I1382 (.Y(inst_cellmath__37[16]), .A(N5562), .B(N5348), .S0(N5360));
INVXL mx2i_A_I4781 (.Y(N10862), .A(N5360));
AOI22XL mx2i_A_I4782 (.Y(inst_cellmath__37[17]), .A0(N5423), .A1(N10862), .B0(N5360), .B1(N5405));
MXI2X2 inst_cellmath__37_0_I1384 (.Y(inst_cellmath__37[18]), .A(N5529), .B(N5458), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1385 (.Y(inst_cellmath__37[19]), .A(N5390), .B(N5511), .S0(N5360));
MXI2X1 inst_cellmath__37_0_I1386 (.Y(inst_cellmath__37[20]), .A(N5445), .B(N5567), .S0(N5360));
MXI2X1 inst_cellmath__37_0_I1387 (.Y(inst_cellmath__37[21]), .A(N5498), .B(N5372), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1388 (.Y(inst_cellmath__37[22]), .A(N5554), .B(N5426), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1389 (.Y(inst_cellmath__37[23]), .A(N5357), .B(N5479), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1390 (.Y(inst_cellmath__37[24]), .A(N5415), .B(N5534), .S0(N5360));
MXI2X1 inst_cellmath__37_0_I1392 (.Y(inst_cellmath__37[26]), .A(N5521), .B(N5394), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1393 (.Y(inst_cellmath__37[27]), .A(N5577), .B(N5501), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1394 (.Y(inst_cellmath__37[28]), .A(N5382), .B(N5362), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1395 (.Y(inst_cellmath__37[29]), .A(N5436), .B(N5470), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1396 (.Y(inst_cellmath__37[30]), .A(N5489), .B(N5579), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1397 (.Y(inst_cellmath__37[31]), .A(N5544), .B(N5440), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1398 (.Y(inst_cellmath__37[32]), .A(N5348), .B(N5547), .S0(N5360));
MXI2XL inst_cellmath__37_0_I1399 (.Y(inst_cellmath__37[33]), .A(N5405), .B(N5407), .S0(N5360));
MXI2XL inst_cellmath__33_49_24_I10972 (.Y(N17372), .A(N5467), .B(N5338), .S0(N5360));
OR2XL inst_cellmath__33_49_24_I11182 (.Y(N17391), .A(inst_cellmath__16), .B(inst_cellmath__11));
NOR2X2 inst_cellmath__33_49_24_I10973 (.Y(N5837), .A(inst_cellmath__30), .B(N17391));
AND2XL inst_cellmath__33_49_24_I10974 (.Y(inst_cellmath__33[24]), .A(N5837), .B(inst_cellmath__37[24]));
NOR2XL inst_cellmath__42__22__I1450 (.Y(N5931), .A(inst_cellmath__37[10]), .B(inst_cellmath__37[23]));
NOR2XL inst_cellmath__42__22__I1449 (.Y(N5919), .A(inst_cellmath__37[11]), .B(inst_cellmath__37[19]));
NOR3X1 inst_cellmath__42__22__I1443 (.Y(N5922), .A(inst_cellmath__30), .B(inst_cellmath__37[2]), .C(inst_cellmath__37[5]));
NOR2X1 inst_cellmath__42__22__I1447 (.Y(N5901), .A(inst_cellmath__37[8]), .B(inst_cellmath__37[16]));
NAND2X2 inst_cellmath__42__22__I1454 (.Y(N5899), .A(N5922), .B(N5901));
OR3XL inst_cellmath__42__22__I1451 (.Y(N5894), .A(inst_cellmath__37[4]), .B(inst_cellmath__37[3]), .C(inst_cellmath__37[22]));
NOR2XL inst_cellmath__42__22__I1445 (.Y(N5926), .A(inst_cellmath__37[9]), .B(inst_cellmath__37[12]));
NOR2X1 inst_cellmath__42__22__I1446 (.Y(N5892), .A(inst_cellmath__37[13]), .B(inst_cellmath__37[14]));
NAND2X1 inst_cellmath__42__22__I1453 (.Y(N5890), .A(N5926), .B(N5892));
OR3X1 inst_cellmath__42__22__I1452 (.Y(N5924), .A(inst_cellmath__37[7]), .B(inst_cellmath__37[15]), .C(inst_cellmath__37[17]));
NOR2X1 inst_cellmath__42__22__I1448 (.Y(N5909), .A(inst_cellmath__37[21]), .B(inst_cellmath__37[20]));
NOR3X1 inst_cellmath__42__22__I1444 (.Y(N5905), .A(inst_cellmath__37[0]), .B(inst_cellmath__37[6]), .C(inst_cellmath__37[1]));
NAND2X2 inst_cellmath__42__22__I1456 (.Y(N5916), .A(N5905), .B(N5909));
CLKAND2X2 inst_cellmath__33_49_24_I11176 (.Y(N17808), .A(N5931), .B(N5919));
NOR2X4 inst_cellmath__33_49_24_I11177 (.Y(N17814), .A(inst_cellmath__37[18]), .B(N5899));
NOR2X2 inst_cellmath__33_49_24_I11178 (.Y(N17821), .A(N5894), .B(N5890));
NOR2X4 inst_cellmath__33_49_24_I11179 (.Y(N17828), .A(N5916), .B(N5924));
NAND2X6 inst_cellmath__33_49_24_I11180 (.Y(N17835), .A(N17814), .B(N17808));
NAND2X4 inst_cellmath__33_49_24_I11181 (.Y(N17811), .A(N17821), .B(N17828));
NOR2XL inst_cellmath__33_49_24_I11183 (.Y(N17829), .A(inst_cellmath__11), .B(inst_cellmath__16));
OAI21X4 inst_cellmath__33_49_24_I11184 (.Y(N17393), .A0(N17835), .A1(N17811), .B0(N17829));
INVXL inst_cellmath__33_49_24_I10977 (.Y(N5967), .A(inst_cellmath__39[25]));
NOR2X2 inst_cellmath__33_49_24_I10978 (.Y(N17379), .A(N5967), .B(inst_cellmath__33[24]));
DLY1X1 inst_cellmath__33_49_24_I10979 (.Y(N5955), .A(N17393));
NAND2XL inst_cellmath__33_49_24_I10980 (.Y(inst_cellmath__44), .A(N17379), .B(N5955));
NAND2XL inst_cellmath__33_49_24_I10981 (.Y(N17371), .A(N5837), .B(N17372));
XOR2XL inst_cellmath__33_49_24_I10982 (.Y(inst_cellmath__39[0]), .A(N17371), .B(inst_cellmath__39[25]));
NAND3BX4 inst_cellmath__33_49_24_I10983 (.Y(N6295), .AN(inst_cellmath__39[0]), .B(N17379), .C(N17393));
AND2XL inst_cellmath__33_49_24_I1420 (.Y(inst_cellmath__33[27]), .A(N5837), .B(inst_cellmath__37[27]));
AND2XL inst_cellmath__33_49_24_I1421 (.Y(inst_cellmath__33[28]), .A(N5837), .B(inst_cellmath__37[28]));
AND2XL inst_cellmath__33_49_24_I1422 (.Y(inst_cellmath__33[29]), .A(N5837), .B(inst_cellmath__37[29]));
AND2XL inst_cellmath__33_49_24_I1424 (.Y(inst_cellmath__33[31]), .A(N5837), .B(inst_cellmath__37[31]));
NAND2XL inst_cellmath__33_49_24_I1426 (.Y(inst_cellmath__33[33]), .A(N5837), .B(inst_cellmath__37[33]));
NOR3BXL inst_cellmath__33_49_24_I4347 (.Y(inst_cellmath__33[34]), .AN(N5837), .B(N5360), .C(N5458));
NOR3BXL inst_cellmath__33_49_24_I4348 (.Y(inst_cellmath__33[35]), .AN(N5837), .B(N5360), .C(N5511));
NOR3BXL inst_cellmath__33_49_24_I4349 (.Y(inst_cellmath__33[36]), .AN(N5837), .B(N5360), .C(N5567));
NOR3BXL inst_cellmath__33_49_24_I4350 (.Y(inst_cellmath__33[37]), .AN(N5837), .B(N5360), .C(N5372));
NOR3BXL inst_cellmath__33_49_24_I4351 (.Y(inst_cellmath__33[38]), .AN(N5837), .B(N5360), .C(N5426));
NOR3BXL inst_cellmath__33_49_24_I4352 (.Y(inst_cellmath__33[39]), .AN(N5837), .B(N5479), .C(N5360));
NOR3BXL inst_cellmath__33_49_24_I4353 (.Y(inst_cellmath__33[40]), .AN(N5837), .B(N5360), .C(N5534));
NOR3BXL inst_cellmath__33_49_24_I4354 (.Y(inst_cellmath__33[41]), .AN(N5837), .B(N5360), .C(N5338));
NOR3BXL inst_cellmath__33_49_24_I4355 (.Y(inst_cellmath__33[42]), .AN(N5837), .B(N5360), .C(N5394));
NOR3BXL inst_cellmath__33_49_24_I4356 (.Y(inst_cellmath__33[43]), .AN(N5837), .B(N5360), .C(N5501));
NOR3BXL inst_cellmath__33_49_24_I4357 (.Y(inst_cellmath__33[44]), .AN(N5837), .B(N5360), .C(N5362));
NOR3BXL inst_cellmath__33_49_24_I4358 (.Y(inst_cellmath__33[45]), .AN(N5837), .B(N5360), .C(N5470));
NOR3BXL inst_cellmath__33_49_24_I4359 (.Y(inst_cellmath__33[46]), .AN(N5837), .B(N5360), .C(N5579));
NOR3BXL inst_cellmath__33_49_24_I4360 (.Y(inst_cellmath__33[47]), .AN(N5837), .B(N5360), .C(N5440));
NOR3BXL inst_cellmath__33_49_24_I4361 (.Y(inst_cellmath__33[48]), .AN(N5837), .B(N5360), .C(N5547));
NOR3BXL inst_cellmath__33_49_24_I4362 (.Y(inst_cellmath__33[49]), .AN(N5837), .B(N5360), .C(N5407));
INVXL cynw_cm_float_add2_ieee_I11281 (.Y(N1693), .A(N5955));
INVXL inst_cellmath__40_I1469 (.Y(N6017), .A(N4309));
INVXL inst_cellmath__40_I1470 (.Y(N6023), .A(N6017));
MX2XL inst_cellmath__40_I1471 (.Y(N655), .A(a_man[0]), .B(b_man[0]), .S0(N6023));
MX2XL inst_cellmath__40_I1472 (.Y(N656), .A(a_man[1]), .B(b_man[1]), .S0(N6023));
MX2XL inst_cellmath__40_I1473 (.Y(N657), .A(a_man[2]), .B(b_man[2]), .S0(N6023));
MX2XL inst_cellmath__40_I1475 (.Y(N658), .A(a_man[3]), .B(b_man[3]), .S0(N6023));
MX2XL inst_cellmath__40_I1476 (.Y(N659), .A(a_man[4]), .B(b_man[4]), .S0(N6023));
MX2XL inst_cellmath__40_I1477 (.Y(N660), .A(a_man[5]), .B(b_man[5]), .S0(N6023));
MX2XL inst_cellmath__40_I1478 (.Y(N661), .A(a_man[6]), .B(b_man[6]), .S0(N6023));
MX2XL inst_cellmath__40_I1479 (.Y(N662), .A(a_man[7]), .B(b_man[7]), .S0(N6023));
MX2XL inst_cellmath__40_I1481 (.Y(N663), .A(a_man[8]), .B(b_man[8]), .S0(N6023));
MX2XL inst_cellmath__40_I1482 (.Y(N664), .A(a_man[9]), .B(b_man[9]), .S0(N6023));
MX2XL inst_cellmath__40_I1483 (.Y(N665), .A(a_man[10]), .B(b_man[10]), .S0(N6023));
MX2XL inst_cellmath__40_I1484 (.Y(N666), .A(a_man[11]), .B(b_man[11]), .S0(N6023));
MX2XL inst_cellmath__40_I1485 (.Y(N667), .A(a_man[12]), .B(b_man[12]), .S0(N6023));
MX2XL inst_cellmath__40_I1487 (.Y(N668), .A(a_man[13]), .B(b_man[13]), .S0(N6023));
MX2XL inst_cellmath__40_I1488 (.Y(N669), .A(a_man[14]), .B(b_man[14]), .S0(N6023));
MX2XL inst_cellmath__40_I1490 (.Y(N671), .A(a_man[16]), .B(b_man[16]), .S0(N6023));
MX2XL inst_cellmath__40_I1491 (.Y(N672), .A(a_man[17]), .B(b_man[17]), .S0(N6023));
MX2XL inst_cellmath__40_I1492 (.Y(N673), .A(a_man[18]), .B(b_man[18]), .S0(N6023));
MX2XL inst_cellmath__40_I1493 (.Y(N674), .A(a_man[19]), .B(b_man[19]), .S0(N6023));
MX2XL inst_cellmath__40_I1494 (.Y(N675), .A(a_man[20]), .B(b_man[20]), .S0(N6023));
MX2XL inst_cellmath__40_I1495 (.Y(N676), .A(a_man[21]), .B(b_man[21]), .S0(N6023));
MX2XL inst_cellmath__40_I1496 (.Y(N677), .A(a_man[22]), .B(b_man[22]), .S0(N6023));
NAND2XL node_cs_const1_cs_ii_A_I4743 (.Y(N10782), .A(N5837), .B(inst_cellmath__37[26]));
CLKXOR2X1 node_cs_const1_cs_ii_A_I4744 (.Y(inst_cellmath__39[1]), .A(N5967), .B(N10782));
XNOR2X1 inst_cellmath__39__19__2mx_I1500 (.Y(inst_cellmath__39[2]), .A(N5967), .B(inst_cellmath__33[27]));
XNOR2X1 inst_cellmath__39__19__2mx_I1501 (.Y(inst_cellmath__39[3]), .A(N5967), .B(inst_cellmath__33[28]));
XNOR2X1 inst_cellmath__39__19__2mx_I1502 (.Y(inst_cellmath__39[4]), .A(N5967), .B(inst_cellmath__33[29]));
NAND2XL node_cs_const1_cs_ii_A_I11454 (.Y(N17952), .A(N5837), .B(inst_cellmath__37[30]));
XOR2XL node_cs_const1_cs_ii_A_I11455 (.Y(inst_cellmath__39[5]), .A(N5967), .B(N17952));
XNOR2X1 inst_cellmath__39__19__2mx_I1504 (.Y(inst_cellmath__39[6]), .A(N5967), .B(inst_cellmath__33[31]));
NAND2XL node_cs_const1_cs_ii_A_I11456 (.Y(N17959), .A(N5837), .B(inst_cellmath__37[32]));
XOR2XL node_cs_const1_cs_ii_A_I11457 (.Y(inst_cellmath__39[7]), .A(N5967), .B(N17959));
CLKXOR2X1 inst_cellmath__39__19__2mx_I4572 (.Y(inst_cellmath__39[8]), .A(N5967), .B(inst_cellmath__33[33]));
XNOR2XL inst_cellmath__39__19__2mx_I1508 (.Y(inst_cellmath__39[9]), .A(N5967), .B(inst_cellmath__33[34]));
XNOR2X1 inst_cellmath__39__19__2mx_I1509 (.Y(inst_cellmath__39[10]), .A(N5967), .B(inst_cellmath__33[35]));
XNOR2X1 inst_cellmath__39__19__2mx_I1510 (.Y(inst_cellmath__39[11]), .A(N5967), .B(inst_cellmath__33[36]));
XNOR2X1 inst_cellmath__39__19__2mx_I1511 (.Y(inst_cellmath__39[12]), .A(N5967), .B(inst_cellmath__33[37]));
XNOR2X1 inst_cellmath__39__19__2mx_I1512 (.Y(inst_cellmath__39[13]), .A(N5967), .B(inst_cellmath__33[38]));
XNOR2X1 inst_cellmath__39__19__2mx_I1513 (.Y(inst_cellmath__39[14]), .A(N5967), .B(inst_cellmath__33[39]));
XNOR2X1 inst_cellmath__39__19__2mx_I1514 (.Y(inst_cellmath__39[15]), .A(N5967), .B(inst_cellmath__33[40]));
XNOR2X1 inst_cellmath__39__19__2mx_I1516 (.Y(inst_cellmath__39[17]), .A(N5967), .B(inst_cellmath__33[42]));
XNOR2X1 inst_cellmath__39__19__2mx_I1517 (.Y(inst_cellmath__39[18]), .A(N5967), .B(inst_cellmath__33[43]));
XNOR2X1 inst_cellmath__39__19__2mx_I1518 (.Y(inst_cellmath__39[19]), .A(N5967), .B(inst_cellmath__33[44]));
XNOR2X1 inst_cellmath__39__19__2mx_I1519 (.Y(inst_cellmath__39[20]), .A(N5967), .B(inst_cellmath__33[45]));
XNOR2X1 inst_cellmath__39__19__2mx_I1520 (.Y(inst_cellmath__39[21]), .A(N5967), .B(inst_cellmath__33[46]));
XNOR2X1 inst_cellmath__39__19__2mx_I1521 (.Y(inst_cellmath__39[22]), .A(N5967), .B(inst_cellmath__33[47]));
XNOR2X1 inst_cellmath__39__19__2mx_I1522 (.Y(inst_cellmath__39[23]), .A(N5967), .B(inst_cellmath__33[48]));
NOR2X2 inst_cellmath__45_0_I1525 (.Y(N6367), .A(inst_cellmath__39[1]), .B(N655));
NAND2X2 inst_cellmath__45_0_I1526 (.Y(N6437), .A(N655), .B(inst_cellmath__39[1]));
NOR2X1 inst_cellmath__45_0_I1527 (.Y(N6179), .A(N656), .B(inst_cellmath__39[2]));
NAND2X1 inst_cellmath__45_0_I1528 (.Y(N6254), .A(N656), .B(inst_cellmath__39[2]));
NOR2XL inst_cellmath__45_0_I1529 (.Y(N6325), .A(N657), .B(inst_cellmath__39[3]));
NAND2X1 inst_cellmath__45_0_I1530 (.Y(N6394), .A(inst_cellmath__39[3]), .B(N657));
NOR2X1 inst_cellmath__45_0_I1531 (.Y(N6467), .A(N658), .B(inst_cellmath__39[4]));
NAND2X2 inst_cellmath__45_0_I1532 (.Y(N6211), .A(N658), .B(inst_cellmath__39[4]));
NOR2XL inst_cellmath__45_0_I1533 (.Y(N6281), .A(N659), .B(inst_cellmath__39[5]));
NAND2X1 inst_cellmath__45_0_I1534 (.Y(N6355), .A(N659), .B(inst_cellmath__39[5]));
NOR2X1 inst_cellmath__45_0_I1535 (.Y(N6424), .A(N660), .B(inst_cellmath__39[6]));
NAND2X1 inst_cellmath__45_0_I1536 (.Y(N6167), .A(N660), .B(inst_cellmath__39[6]));
NOR2XL inst_cellmath__45_0_I1537 (.Y(N6240), .A(N661), .B(inst_cellmath__39[7]));
NAND2X1 inst_cellmath__45_0_I1538 (.Y(N6312), .A(N661), .B(inst_cellmath__39[7]));
NOR2X1 inst_cellmath__45_0_I1539 (.Y(N6381), .A(N662), .B(inst_cellmath__39[8]));
NAND2X2 inst_cellmath__45_0_I1540 (.Y(N6452), .A(N662), .B(inst_cellmath__39[8]));
NOR2XL inst_cellmath__45_0_I1541 (.Y(N6195), .A(N663), .B(inst_cellmath__39[9]));
NAND2XL inst_cellmath__45_0_I1542 (.Y(N6268), .A(N663), .B(inst_cellmath__39[9]));
NOR2XL inst_cellmath__45_0_I1543 (.Y(N6342), .A(N664), .B(inst_cellmath__39[10]));
NAND2XL inst_cellmath__45_0_I1544 (.Y(N6411), .A(N664), .B(inst_cellmath__39[10]));
NOR2XL inst_cellmath__45_0_I1545 (.Y(N6156), .A(N665), .B(inst_cellmath__39[11]));
NAND2XL inst_cellmath__45_0_I1546 (.Y(N6229), .A(N665), .B(inst_cellmath__39[11]));
NOR2XL inst_cellmath__45_0_I1547 (.Y(N6302), .A(N666), .B(inst_cellmath__39[12]));
NAND2XL inst_cellmath__45_0_I1548 (.Y(N6373), .A(N666), .B(inst_cellmath__39[12]));
NOR2XL inst_cellmath__45_0_I1549 (.Y(N6443), .A(N667), .B(inst_cellmath__39[13]));
NAND2XL inst_cellmath__45_0_I1550 (.Y(N6185), .A(N667), .B(inst_cellmath__39[13]));
NOR2XL inst_cellmath__45_0_I1551 (.Y(N6261), .A(N668), .B(inst_cellmath__39[14]));
NAND2XL inst_cellmath__45_0_I1552 (.Y(N6331), .A(N668), .B(inst_cellmath__39[14]));
NOR2XL inst_cellmath__45_0_I1553 (.Y(N6401), .A(N669), .B(inst_cellmath__39[15]));
NAND2XL inst_cellmath__45_0_I1554 (.Y(N6473), .A(N669), .B(inst_cellmath__39[15]));
NOR2XL inst_cellmath__45_0_I1557 (.Y(N6362), .A(N671), .B(inst_cellmath__39[17]));
NAND2XL inst_cellmath__45_0_I1558 (.Y(N6430), .A(N671), .B(inst_cellmath__39[17]));
NOR2XL inst_cellmath__45_0_I1559 (.Y(N6173), .A(N672), .B(inst_cellmath__39[18]));
NAND2XL inst_cellmath__45_0_I1560 (.Y(N6247), .A(N672), .B(inst_cellmath__39[18]));
NOR2XL inst_cellmath__45_0_I1561 (.Y(N6318), .A(N673), .B(inst_cellmath__39[19]));
NAND2XL inst_cellmath__45_0_I1562 (.Y(N6388), .A(N673), .B(inst_cellmath__39[19]));
NOR2XL inst_cellmath__45_0_I1563 (.Y(N6460), .A(N674), .B(inst_cellmath__39[20]));
NAND2XL inst_cellmath__45_0_I1564 (.Y(N6202), .A(N674), .B(inst_cellmath__39[20]));
NOR2XL inst_cellmath__45_0_I1565 (.Y(N6274), .A(N675), .B(inst_cellmath__39[21]));
NAND2XL inst_cellmath__45_0_I1566 (.Y(N6347), .A(N675), .B(inst_cellmath__39[21]));
NOR2XL inst_cellmath__45_0_I1567 (.Y(N6416), .A(N676), .B(inst_cellmath__39[22]));
NAND2XL inst_cellmath__45_0_I1568 (.Y(N6161), .A(N676), .B(inst_cellmath__39[22]));
NOR2XL inst_cellmath__45_0_I1569 (.Y(N6233), .A(N677), .B(inst_cellmath__39[23]));
NAND2XL inst_cellmath__45_0_I1570 (.Y(N6305), .A(N677), .B(inst_cellmath__39[23]));
XOR2XL inst_cellmath__45_0_I4573 (.Y(N6376), .A(N5967), .B(inst_cellmath__33[49]));
INVXL inst_cellmath__45_0_I1572 (.Y(N6387), .A(N6295));
AOI21X1 inst_cellmath__45_0_I1574 (.Y(N6477), .A0(N6367), .A1(N6254), .B0(N6179));
NAND2XL inst_cellmath__45_0_I1575 (.Y(N6222), .A(N6254), .B(N6437));
AOI21X1 inst_cellmath__45_0_I1578 (.Y(N6435), .A0(N6211), .A1(N6325), .B0(N6467));
NAND2XL inst_cellmath__45_0_I1579 (.Y(N6177), .A(N6394), .B(N6211));
AOI21X1 inst_cellmath__45_0_I1582 (.Y(N6392), .A0(N6167), .A1(N6281), .B0(N6424));
NAND2XL inst_cellmath__45_0_I1583 (.Y(N6465), .A(N6167), .B(N6355));
AOI21X1 inst_cellmath__45_0_I1586 (.Y(N6353), .A0(N6240), .A1(N6452), .B0(N6381));
NAND2XL inst_cellmath__45_0_I1587 (.Y(N6422), .A(N6452), .B(N6312));
AOI21X1 inst_cellmath__45_0_I1588 (.Y(N6165), .A0(N6268), .A1(N6381), .B0(N6195));
NAND2XL inst_cellmath__45_0_I1589 (.Y(N6238), .A(N6268), .B(N6452));
AOI21XL inst_cellmath__45_0_I1590 (.Y(N6310), .A0(N6411), .A1(N6195), .B0(N6342));
NAND2XL inst_cellmath__45_0_I1591 (.Y(N6380), .A(N6411), .B(N6268));
AOI21XL inst_cellmath__45_0_I1592 (.Y(N6451), .A0(N6229), .A1(N6342), .B0(N6156));
NAND2XL inst_cellmath__45_0_I1593 (.Y(N6194), .A(N6229), .B(N6411));
AOI21XL inst_cellmath__45_0_I1594 (.Y(N6267), .A0(N6373), .A1(N6156), .B0(N6302));
NAND2XL inst_cellmath__45_0_I1595 (.Y(N6341), .A(N6373), .B(N6229));
AOI21XL inst_cellmath__45_0_I1596 (.Y(N6410), .A0(N6185), .A1(N6302), .B0(N6443));
NAND2XL inst_cellmath__45_0_I1597 (.Y(N6155), .A(N6185), .B(N6373));
AOI21XL inst_cellmath__45_0_I1598 (.Y(N6228), .A0(N6331), .A1(N6443), .B0(N6261));
NAND2XL inst_cellmath__45_0_I1599 (.Y(N6300), .A(N6331), .B(N6185));
AOI21XL inst_cellmath__45_0_I1600 (.Y(N6372), .A0(N6473), .A1(N6261), .B0(N6401));
NAND2XL inst_cellmath__45_0_I1601 (.Y(N6442), .A(N6473), .B(N6331));
MX2XL inst_cellmath__45_0_I11149 (.Y(N17769), .A(a_man[15]), .B(b_man[15]), .S0(N6023));
XNOR2X1 inst_cellmath__45_0_I11150 (.Y(N17778), .A(N5967), .B(inst_cellmath__33[41]));
NAND2XL inst_cellmath__45_0_I11152 (.Y(N6287), .A(N17769), .B(N17778));
NOR2XL inst_cellmath__45_0_I11151 (.Y(N6218), .A(N17769), .B(N17778));
AOI21XL inst_cellmath__45_0_I1602 (.Y(N6184), .A0(N6287), .A1(N6401), .B0(N6218));
NAND2XL inst_cellmath__45_0_I1603 (.Y(N6260), .A(N6287), .B(N6473));
AOI21XL inst_cellmath__45_0_I1604 (.Y(N6330), .A0(N6430), .A1(N6218), .B0(N6362));
NAND2XL inst_cellmath__45_0_I1605 (.Y(N6400), .A(N6430), .B(N6287));
AOI21XL inst_cellmath__45_0_I1606 (.Y(N6472), .A0(N6247), .A1(N6362), .B0(N6173));
NAND2XL inst_cellmath__45_0_I1607 (.Y(N6217), .A(N6247), .B(N6430));
AOI21XL inst_cellmath__45_0_I1608 (.Y(N6286), .A0(N6388), .A1(N6173), .B0(N6318));
NAND2XL inst_cellmath__45_0_I1609 (.Y(N6360), .A(N6388), .B(N6247));
AOI21XL inst_cellmath__45_0_I1610 (.Y(N6429), .A0(N6202), .A1(N6318), .B0(N6460));
NAND2XL inst_cellmath__45_0_I1611 (.Y(N6172), .A(N6202), .B(N6388));
AOI21XL inst_cellmath__45_0_I1612 (.Y(N6245), .A0(N6347), .A1(N6460), .B0(N6274));
NAND2XL inst_cellmath__45_0_I1613 (.Y(N6317), .A(N6347), .B(N6202));
AOI21XL inst_cellmath__45_0_I1614 (.Y(N6386), .A0(N6161), .A1(N6274), .B0(N6416));
NAND2XL inst_cellmath__45_0_I1615 (.Y(N6457), .A(N6161), .B(N6347));
AOI21XL inst_cellmath__45_0_I1616 (.Y(N6200), .A0(N6305), .A1(N6416), .B0(N6233));
NAND2XL inst_cellmath__45_0_I1617 (.Y(N6272), .A(N6305), .B(N6161));
NAND2XL inst_cellmath__45_0_I1618 (.Y(N6159), .A(N6376), .B(N6305));
INVXL inst_cellmath__45_0_I1619 (.Y(N6459), .A(N6387));
AOI21X2 inst_cellmath__45_0_I11094 (.Y(N6336), .A0(N6437), .A1(N6295), .B0(N6367));
INVXL inst_cellmath__45_0_I1620 (.Y(N6201), .A(N6336));
OAI21X1 inst_cellmath__45_0_I1621 (.Y(N6475), .A0(N6222), .A1(N6387), .B0(N6477));
OAI21X1 inst_cellmath__45_0_I1623 (.Y(N6432), .A0(N6177), .A1(N6477), .B0(N6435));
NOR2X1 inst_cellmath__45_0_I1624 (.Y(N6176), .A(N6177), .B(N6222));
NAND2XL inst_cellmath__45_0_I11098 (.Y(N6323), .A(N6355), .B(N6211));
AOI21X1 inst_cellmath__45_0_I11095 (.Y(N6293), .A0(N6179), .A1(N6394), .B0(N6325));
AOI21XL inst_cellmath__45_0_I11097 (.Y(N6252), .A0(N6467), .A1(N6355), .B0(N6281));
OAI21XL inst_cellmath__45_0_I1625 (.Y(N6250), .A0(N6323), .A1(N6293), .B0(N6252));
NAND2XL inst_cellmath__45_0_I11096 (.Y(N6365), .A(N6254), .B(N6394));
NOR2X1 inst_cellmath__45_0_I1626 (.Y(N6321), .A(N6365), .B(N6323));
OAI21XL inst_cellmath__45_0_I1627 (.Y(N6390), .A0(N6465), .A1(N6435), .B0(N6392));
NOR2XL inst_cellmath__45_0_I1628 (.Y(N6463), .A(N6465), .B(N6177));
OAI21XL inst_cellmath__45_0_I1631 (.Y(N6350), .A0(N6422), .A1(N6392), .B0(N6353));
NOR2XL inst_cellmath__45_0_I1632 (.Y(N6419), .A(N6422), .B(N6465));
AOI21XL inst_cellmath__45_0_I11099 (.Y(N6209), .A0(N6424), .A1(N6312), .B0(N6240));
OAI21XL inst_cellmath__45_0_I1633 (.Y(N6164), .A0(N6238), .A1(N6209), .B0(N6165));
NAND2XL inst_cellmath__45_0_I11100 (.Y(N6279), .A(N6167), .B(N6312));
NOR2XL inst_cellmath__45_0_I1634 (.Y(N6236), .A(N6238), .B(N6279));
OAI21X1 inst_cellmath__45_0_I1635 (.Y(N6308), .A0(N6380), .A1(N6353), .B0(N6310));
NOR2XL inst_cellmath__45_0_I1636 (.Y(N6379), .A(N6380), .B(N6422));
OAI21XL inst_cellmath__45_0_I1639 (.Y(N6266), .A0(N6341), .A1(N6310), .B0(N6267));
NOR2XL inst_cellmath__45_0_I1640 (.Y(N6340), .A(N6341), .B(N6380));
OAI21XL inst_cellmath__45_0_I1641 (.Y(N6408), .A0(N6155), .A1(N6451), .B0(N6410));
NOR2XL inst_cellmath__45_0_I1642 (.Y(N6154), .A(N6155), .B(N6194));
OAI21XL inst_cellmath__45_0_I1643 (.Y(N6227), .A0(N6300), .A1(N6267), .B0(N6228));
NOR2XL inst_cellmath__45_0_I1644 (.Y(N6298), .A(N6300), .B(N6341));
OAI21XL inst_cellmath__45_0_I1647 (.Y(N6182), .A0(N6260), .A1(N6228), .B0(N6184));
NOR2XL inst_cellmath__45_0_I1648 (.Y(N6258), .A(N6260), .B(N6300));
OAI21XL inst_cellmath__45_0_I1649 (.Y(N6329), .A0(N6400), .A1(N6372), .B0(N6330));
NOR2XL inst_cellmath__45_0_I1650 (.Y(N6397), .A(N6400), .B(N6442));
OAI21XL inst_cellmath__45_0_I1651 (.Y(N6471), .A0(N6217), .A1(N6184), .B0(N6472));
NOR2XL inst_cellmath__45_0_I1652 (.Y(N6215), .A(N6217), .B(N6260));
OAI21XL inst_cellmath__45_0_I1653 (.Y(N6284), .A0(N6360), .A1(N6330), .B0(N6286));
NOR2XL inst_cellmath__45_0_I1654 (.Y(N6359), .A(N6360), .B(N6400));
OAI21XL inst_cellmath__45_0_I1655 (.Y(N6428), .A0(N6172), .A1(N6472), .B0(N6429));
NOR2XL inst_cellmath__45_0_I1656 (.Y(N6170), .A(N6172), .B(N6217));
OAI21XL inst_cellmath__45_0_I1657 (.Y(N6244), .A0(N6317), .A1(N6286), .B0(N6245));
NOR2XL inst_cellmath__45_0_I1658 (.Y(N6316), .A(N6317), .B(N6360));
OAI21XL inst_cellmath__45_0_I1659 (.Y(N6384), .A0(N6457), .A1(N6429), .B0(N6386));
NOR2XL inst_cellmath__45_0_I1660 (.Y(N6456), .A(N6457), .B(N6172));
OAI21XL inst_cellmath__45_0_I1661 (.Y(N6199), .A0(N6272), .A1(N6245), .B0(N6200));
NOR2XL inst_cellmath__45_0_I1662 (.Y(N6270), .A(N6272), .B(N6317));
OAI2BB2XL inst_cellmath__45_0_I1663 (.Y(N6344), .A0N(N6376), .A1N(N6233), .B0(N6159), .B1(N6386));
NOR2XL inst_cellmath__45_0_I1664 (.Y(N6413), .A(N6159), .B(N6457));
INVXL inst_cellmath__45_0_I1665 (.Y(N6273), .A(N6459));
INVXL inst_cellmath__45_0_I1666 (.Y(N6346), .A(N6201));
INVXL inst_cellmath__45_0_I1667 (.Y(N6415), .A(N6475));
OAI21X2 inst_cellmath__45_0_I11160 (.Y(N6291), .A0(N6365), .A1(N6336), .B0(N6293));
INVXL inst_cellmath__45_0_I1668 (.Y(N6160), .A(N6291));
AOI21XL inst_cellmath__45_0_I1669 (.Y(N6220), .A0(N6176), .A1(N6459), .B0(N6432));
AOI21X1 inst_cellmath__45_0_I1670 (.Y(N6363), .A0(N6321), .A1(N6201), .B0(N6250));
AOI21X1 inst_cellmath__45_0_I1671 (.Y(N6174), .A0(N6463), .A1(N6475), .B0(N6390));
AOI21X1 inst_cellmath__45_0_I1673 (.Y(N6461), .A0(N6419), .A1(N6432), .B0(N6350));
NAND2XL inst_cellmath__45_0_I1674 (.Y(N6204), .A(N6176), .B(N6419));
AOI21X1 inst_cellmath__45_0_I1675 (.Y(N6275), .A0(N6236), .A1(N6250), .B0(N6164));
NAND2XL inst_cellmath__45_0_I1676 (.Y(N6348), .A(N6236), .B(N6321));
AOI21X1 inst_cellmath__45_0_I1677 (.Y(N6418), .A0(N6379), .A1(N6390), .B0(N6308));
NAND2XL inst_cellmath__45_0_I1678 (.Y(N6162), .A(N6379), .B(N6463));
NOR2X1 inst_cellmath__45_0_I11154 (.Y(N6192), .A(N6238), .B(N6194));
OAI21X1 inst_cellmath__45_0_I11161 (.Y(N6205), .A0(N6279), .A1(N6252), .B0(N6209));
OAI21X1 inst_cellmath__45_0_I11153 (.Y(N6450), .A0(N6194), .A1(N6165), .B0(N6451));
AOI21X1 inst_cellmath__45_0_I1679 (.Y(N6234), .A0(N6192), .A1(N6205), .B0(N6450));
NOR2XL inst_cellmath__45_0_I11159 (.Y(N6277), .A(N6323), .B(N6279));
NAND2XL inst_cellmath__45_0_I1680 (.Y(N6307), .A(N6192), .B(N6277));
AOI21XL inst_cellmath__45_0_I1681 (.Y(N6377), .A0(N6340), .A1(N6350), .B0(N6266));
NAND2XL inst_cellmath__45_0_I1682 (.Y(N6448), .A(N6340), .B(N6419));
AOI21X1 inst_cellmath__45_0_I1683 (.Y(N6191), .A0(N6154), .A1(N6164), .B0(N6408));
NAND2XL inst_cellmath__45_0_I1684 (.Y(N6264), .A(N6154), .B(N6236));
AOI21X1 inst_cellmath__45_0_I1685 (.Y(N6338), .A0(N6298), .A1(N6308), .B0(N6227));
NAND2XL inst_cellmath__45_0_I1686 (.Y(N6406), .A(N6379), .B(N6298));
AOI21XL inst_cellmath__45_0_I1689 (.Y(N6296), .A0(N6258), .A1(N6266), .B0(N6182));
NAND2XL inst_cellmath__45_0_I1690 (.Y(N6369), .A(N6258), .B(N6340));
AOI21XL inst_cellmath__45_0_I1691 (.Y(N6439), .A0(N6397), .A1(N6408), .B0(N6329));
NAND2XL inst_cellmath__45_0_I1692 (.Y(N6180), .A(N6397), .B(N6154));
AOI21XL inst_cellmath__45_0_I1693 (.Y(N6256), .A0(N6215), .A1(N6227), .B0(N6471));
NAND2XL inst_cellmath__45_0_I1694 (.Y(N6327), .A(N6215), .B(N6298));
OAI21XL inst_cellmath__45_0_I11155 (.Y(N6371), .A0(N6442), .A1(N6410), .B0(N6372));
AOI21XL inst_cellmath__45_0_I1695 (.Y(N6395), .A0(N6359), .A1(N6371), .B0(N6284));
NOR2X1 inst_cellmath__45_0_I11156 (.Y(N6441), .A(N6442), .B(N6155));
NAND2XL inst_cellmath__45_0_I1696 (.Y(N6469), .A(N6359), .B(N6441));
AOI21XL inst_cellmath__45_0_I1697 (.Y(N6213), .A0(N6170), .A1(N6182), .B0(N6428));
NAND2XL inst_cellmath__45_0_I1698 (.Y(N6282), .A(N6170), .B(N6258));
AOI21XL inst_cellmath__45_0_I1699 (.Y(N6357), .A0(N6316), .A1(N6329), .B0(N6244));
NAND2XL inst_cellmath__45_0_I1700 (.Y(N6426), .A(N6316), .B(N6397));
AOI21XL inst_cellmath__45_0_I1701 (.Y(N6168), .A0(N6456), .A1(N6471), .B0(N6384));
NAND2XL inst_cellmath__45_0_I1702 (.Y(N6242), .A(N6456), .B(N6215));
AOI21XL inst_cellmath__45_0_I1703 (.Y(N6314), .A0(N6270), .A1(N6284), .B0(N6199));
NAND2XL inst_cellmath__45_0_I1704 (.Y(N6382), .A(N6270), .B(N6359));
AOI21XL inst_cellmath__45_0_I1705 (.Y(N6454), .A0(N6413), .A1(N6428), .B0(N6344));
NAND2XL inst_cellmath__45_0_I1706 (.Y(N6197), .A(N6413), .B(N6170));
INVXL inst_cellmath__45_0_I1707 (.Y(N6232), .A(N6273));
INVXL inst_cellmath__45_0_I1708 (.Y(N6304), .A(N6346));
INVX1 inst_cellmath__45_0_I1709 (.Y(N6375), .A(N6415));
INVXL inst_cellmath__45_0_I1710 (.Y(N6446), .A(N6160));
INVXL inst_cellmath__45_0_I1711 (.Y(N6189), .A(N6220));
INVX1 inst_cellmath__45_0_I1712 (.Y(N6263), .A(N6363));
INVX1 inst_cellmath__45_0_I1713 (.Y(N6335), .A(N6174));
AOI21X1 inst_cellmath__45_0_I11157 (.Y(N6480), .A0(N6441), .A1(N6450), .B0(N6371));
NAND2X1 inst_cellmath__45_0_I11158 (.Y(N6225), .A(N6441), .B(N6192));
AOI21X2 inst_cellmath__45_0_I11162 (.Y(N6320), .A0(N6277), .A1(N6291), .B0(N6205));
NOR2X1 inst_cellmath__45_0_I11163 (.Y(N17752), .A(N6225), .B(N6320));
OA21X1 inst_cellmath__45_0_I11164 (.Y(N17776), .A0(N6225), .A1(N6320), .B0(N6480));
NAND2BXL inst_cellmath__45_0_I11165 (.Y(N17746), .AN(N6218), .B(N6287));
INVXL inst_cellmath__45_0_I11166 (.Y(N17754), .A(N17776));
NOR2BX2 inst_cellmath__45_0_I11167 (.Y(N17767), .AN(N6480), .B(N17752));
MXI2X1 inst_cellmath__45_0_I11168 (.Y(inst_cellmath__45[16]), .A(N17767), .B(N17754), .S0(N17746));
INVX1 inst_cellmath__45_0_I11105 (.Y(N6403), .A(N6320));
OAI21X1 inst_cellmath__45_0_I1715 (.Y(N6248), .A0(N6204), .A1(N6273), .B0(N6461));
OAI21XL inst_cellmath__45_0_I1716 (.Y(N6447), .A0(N6406), .A1(N6174), .B0(N6338));
OAI21XL inst_cellmath__45_0_I1717 (.Y(N6404), .A0(N6369), .A1(N6461), .B0(N6296));
NOR2XL inst_cellmath__45_0_I1718 (.Y(N6478), .A(N6369), .B(N6204));
OAI21XL inst_cellmath__45_0_I1719 (.Y(N6223), .A0(N6180), .A1(N6275), .B0(N6439));
NOR2XL inst_cellmath__45_0_I1720 (.Y(N6294), .A(N6180), .B(N6348));
OAI21XL inst_cellmath__45_0_I1721 (.Y(N6366), .A0(N6327), .A1(N6418), .B0(N6256));
NOR2X1 inst_cellmath__45_0_I1722 (.Y(N6436), .A(N6327), .B(N6162));
OAI21X1 inst_cellmath__45_0_I1723 (.Y(N6178), .A0(N6469), .A1(N6234), .B0(N6395));
NOR2XL inst_cellmath__45_0_I1724 (.Y(N6253), .A(N6469), .B(N6307));
OAI21XL inst_cellmath__45_0_I1725 (.Y(N6324), .A0(N6282), .A1(N6377), .B0(N6213));
NOR2XL inst_cellmath__45_0_I1726 (.Y(N6393), .A(N6282), .B(N6448));
OAI21X1 inst_cellmath__45_0_I1727 (.Y(N6466), .A0(N6426), .A1(N6191), .B0(N6357));
NOR2XL inst_cellmath__45_0_I1728 (.Y(N6210), .A(N6264), .B(N6426));
OAI21X1 inst_cellmath__45_0_I1729 (.Y(N6280), .A0(N6242), .A1(N6338), .B0(N6168));
NOR2XL inst_cellmath__45_0_I1730 (.Y(N6354), .A(N6406), .B(N6242));
OAI21X1 inst_cellmath__45_0_I1731 (.Y(N6423), .A0(N6382), .A1(N6480), .B0(N6314));
NOR2XL inst_cellmath__45_0_I1732 (.Y(N6166), .A(N6225), .B(N6382));
OAI21XL inst_cellmath__45_0_I1733 (.Y(N6239), .A0(N6197), .A1(N6296), .B0(N6454));
NOR2XL inst_cellmath__45_0_I1734 (.Y(N6311), .A(N6197), .B(N6369));
OA21XL inst_cellmath__45_0_I1735 (.Y(N6464), .A0(N6348), .A1(N6346), .B0(N6275));
OA21XL inst_cellmath__45_0_I1736 (.Y(N6208), .A0(N6162), .A1(N6415), .B0(N6418));
OA21XL inst_cellmath__45_0_I1737 (.Y(N6278), .A0(N6307), .A1(N6160), .B0(N6234));
OA21X1 inst_cellmath__45_0_I1738 (.Y(N6351), .A0(N6448), .A1(N6220), .B0(N6377));
OA21XL inst_cellmath__45_0_I1739 (.Y(N6421), .A0(N6264), .A1(N6363), .B0(N6191));
AOI21X1 inst_cellmath__45_0_I1741 (.Y(N6188), .A0(N6478), .A1(N6232), .B0(N6404));
AOI21X1 inst_cellmath__45_0_I1742 (.Y(N6334), .A0(N6294), .A1(N6304), .B0(N6223));
AOI21X1 inst_cellmath__45_0_I1743 (.Y(N6476), .A0(N6436), .A1(N6375), .B0(N6366));
AOI21X1 inst_cellmath__45_0_I1744 (.Y(N6292), .A0(N6253), .A1(N6446), .B0(N6178));
AOI21X1 inst_cellmath__45_0_I1745 (.Y(N6434), .A0(N6393), .A1(N6189), .B0(N6324));
AOI21X1 inst_cellmath__45_0_I1746 (.Y(N6251), .A0(N6210), .A1(N6263), .B0(N6466));
AOI21X1 inst_cellmath__45_0_I1747 (.Y(N6391), .A0(N6354), .A1(N6335), .B0(N6280));
AOI21X1 inst_cellmath__45_0_I1748 (.Y(N6207), .A0(N6166), .A1(N6403), .B0(N6423));
AOI21X1 inst_cellmath__45_0_I1749 (.Y(N6352), .A0(N6311), .A1(N6248), .B0(N6239));
NAND2BXL inst_cellmath__45_0_I1750 (.Y(N6158), .AN(N6367), .B(N6437));
NAND2BXL inst_cellmath__45_0_I1751 (.Y(N6374), .AN(N6179), .B(N6254));
NAND2BXL inst_cellmath__45_0_I1752 (.Y(N6262), .AN(N6325), .B(N6394));
NAND2BXL inst_cellmath__45_0_I1753 (.Y(N6474), .AN(N6467), .B(N6211));
NAND2BXL inst_cellmath__45_0_I1754 (.Y(N6364), .AN(N6281), .B(N6355));
NAND2BXL inst_cellmath__45_0_I1755 (.Y(N6249), .AN(N6424), .B(N6167));
NAND2BXL inst_cellmath__45_0_I1756 (.Y(N6462), .AN(N6240), .B(N6312));
NAND2BXL inst_cellmath__45_0_I1757 (.Y(N6349), .AN(N6381), .B(N6452));
NAND2BXL inst_cellmath__45_0_I1758 (.Y(N6235), .AN(N6195), .B(N6268));
NAND2BXL inst_cellmath__45_0_I1759 (.Y(N6449), .AN(N6342), .B(N6411));
NAND2BXL inst_cellmath__45_0_I1760 (.Y(N6339), .AN(N6156), .B(N6229));
NAND2BXL inst_cellmath__45_0_I1761 (.Y(N6226), .AN(N6302), .B(N6373));
NAND2BXL inst_cellmath__45_0_I1762 (.Y(N6440), .AN(N6443), .B(N6185));
NAND2BXL inst_cellmath__45_0_I1763 (.Y(N6328), .AN(N6261), .B(N6331));
NAND2BXL inst_cellmath__45_0_I1764 (.Y(N6214), .AN(N6401), .B(N6473));
NAND2BXL inst_cellmath__45_0_I1766 (.Y(N6315), .AN(N6362), .B(N6430));
NAND2BXL inst_cellmath__45_0_I1767 (.Y(N6198), .AN(N6173), .B(N6247));
NAND2BXL inst_cellmath__45_0_I1768 (.Y(N6412), .AN(N6318), .B(N6388));
NAND2BXL inst_cellmath__45_0_I1769 (.Y(N6303), .AN(N6460), .B(N6202));
NAND2BXL inst_cellmath__45_0_I1770 (.Y(N6186), .AN(N6274), .B(N6347));
NAND2BXL inst_cellmath__45_0_I1771 (.Y(N6402), .AN(N6416), .B(N6161));
NAND2BXL inst_cellmath__45_0_I1772 (.Y(N6288), .AN(N6233), .B(N6305));
XOR2XL inst_cellmath__45_0_I1773 (.Y(inst_cellmath__45[0]), .A(inst_cellmath__39[0]), .B(inst_cellmath__44));
XOR2XL inst_cellmath__45_0_I1775 (.Y(inst_cellmath__45[2]), .A(N6374), .B(N6304));
XOR2XL inst_cellmath__45_0_I1776 (.Y(inst_cellmath__45[3]), .A(N6262), .B(N6375));
CLKXOR2X1 inst_cellmath__45_0_I1777 (.Y(inst_cellmath__45[4]), .A(N6446), .B(N6474));
CLKXOR2X1 inst_cellmath__45_0_I1779 (.Y(inst_cellmath__45[6]), .A(N6263), .B(N6249));
XOR2X1 inst_cellmath__45_0_I1780 (.Y(inst_cellmath__45[7]), .A(N6335), .B(N6462));
CLKXOR2X1 inst_cellmath__45_0_I1781 (.Y(inst_cellmath__45[8]), .A(N6403), .B(N6349));
XNOR2X1 inst_cellmath__45_0_I1783 (.Y(inst_cellmath__45[10]), .A(N6464), .B(N6449));
XNOR2X1 inst_cellmath__45_0_I1784 (.Y(inst_cellmath__45[11]), .A(N6339), .B(N6208));
INVXL inst_cellmath__45_0_I1785 (.Y(N6414), .A(N6278));
MXI2X1 inst_cellmath__45_0_I1786 (.Y(inst_cellmath__45[12]), .A(N6278), .B(N6414), .S0(N6226));
INVXL inst_cellmath__45_0_I1788 (.Y(N6187), .A(N6421));
MXI2X1 inst_cellmath__45_0_I1789 (.Y(inst_cellmath__45[14]), .A(N6421), .B(N6187), .S0(N6328));
CLKXOR2X1 inst_cellmath__45_0_I1790 (.Y(inst_cellmath__45[15]), .A(N6214), .B(N6447));
XNOR2X1 inst_cellmath__45_0_I10985 (.Y(inst_cellmath__45[18]), .A(N6198), .B(N6334));
XNOR2X1 inst_cellmath__45_0_I10986 (.Y(inst_cellmath__45[19]), .A(N6412), .B(N6476));
XNOR2X1 inst_cellmath__45_0_I10987 (.Y(inst_cellmath__45[20]), .A(N6303), .B(N6292));
XNOR2X1 inst_cellmath__45_0_I10988 (.Y(inst_cellmath__45[21]), .A(N6186), .B(N6434));
XNOR2X1 inst_cellmath__45_0_I10989 (.Y(inst_cellmath__45[23]), .A(N6288), .B(N6391));
CLKXOR2X1 inst_cellmath__45_0_I10990 (.Y(inst_cellmath__45[25]), .A(inst_cellmath__39[25]), .B(N6352));
NOR2X4 inst_cellmath__45_0_I10991 (.Y(N6795), .A(inst_cellmath__45[19]), .B(inst_cellmath__45[18]));
NOR2X2 inst_cellmath__45_0_I10992 (.Y(N6816), .A(inst_cellmath__45[21]), .B(inst_cellmath__45[20]));
XNOR2X1 inst_cellmath__45_0_I10993 (.Y(inst_cellmath__45[22]), .A(N6402), .B(N6251));
NOR2X2 inst_cellmath__45_0_I10994 (.Y(N6823), .A(inst_cellmath__45[22]), .B(inst_cellmath__45[23]));
XNOR2XL inst_cellmath__45_0_I4440 (.Y(N10745), .A(N6376), .B(N6207));
INVX2 inst_cellmath__45_0_I10995 (.Y(inst_cellmath__45[24]), .A(N10745));
NOR2X4 inst_cellmath__45_0_I10996 (.Y(N6845), .A(inst_cellmath__45[24]), .B(inst_cellmath__45[25]));
NAND2X6 inst_cellmath__45_0_I10997 (.Y(N6773), .A(N6795), .B(N6816));
NAND2X6 inst_cellmath__45_0_I10998 (.Y(N6793), .A(N6823), .B(N6845));
NOR2X6 inst_cellmath__45_0_I10999 (.Y(N6830), .A(N6773), .B(N6793));
XOR2XL inst_cellmath__50_0_I11056 (.Y(inst_cellmath__45[1]), .A(N6232), .B(N6158));
NOR2XL inst_cellmath__49_0_I1802 (.Y(N6763), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[0]));
NOR2BX1 inst_cellmath__49_0_I1803 (.Y(N6807), .AN(inst_cellmath__45[2]), .B(inst_cellmath__45[3]));
CLKXOR2X1 inst_cellmath__50_0_I11057 (.Y(inst_cellmath__45[5]), .A(N6189), .B(N6364));
INVXL inst_cellmath__49_0_I1804 (.Y(N6826), .A(inst_cellmath__45[5]));
OAI21XL inst_cellmath__49_0_I1805 (.Y(N6848), .A0(inst_cellmath__45[4]), .A1(N6807), .B0(N6826));
NOR2X1 inst_cellmath__49_0_I1806 (.Y(N6774), .A(inst_cellmath__45[2]), .B(inst_cellmath__45[3]));
NOR2X2 inst_cellmath__49_0_I1807 (.Y(N6794), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[4]));
NOR2BX1 inst_cellmath__49_0_I1808 (.Y(N6836), .AN(inst_cellmath__45[6]), .B(inst_cellmath__45[7]));
CLKXOR2X1 inst_cellmath__50_0_I11058 (.Y(inst_cellmath__45[9]), .A(N6235), .B(N6248));
INVXL inst_cellmath__49_0_I1809 (.Y(N6856), .A(inst_cellmath__45[9]));
OAI21XL inst_cellmath__49_0_I1810 (.Y(N6783), .A0(inst_cellmath__45[8]), .A1(N6836), .B0(N6856));
NOR2X2 inst_cellmath__49_0_I1811 (.Y(N6802), .A(inst_cellmath__45[6]), .B(inst_cellmath__45[7]));
NOR2X2 inst_cellmath__49_0_I1812 (.Y(N6821), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[8]));
NOR2BX1 inst_cellmath__49_0_I1813 (.Y(N6769), .AN(inst_cellmath__45[10]), .B(inst_cellmath__45[11]));
XNOR2X1 inst_cellmath__50_0_I11059 (.Y(inst_cellmath__45[13]), .A(N6440), .B(N6351));
INVXL inst_cellmath__49_0_I1814 (.Y(N6790), .A(inst_cellmath__45[13]));
OAI21XL inst_cellmath__49_0_I1815 (.Y(N6812), .A0(inst_cellmath__45[12]), .A1(N6769), .B0(N6790));
NOR2X2 inst_cellmath__49_0_I1816 (.Y(N6832), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[10]));
NOR2X2 inst_cellmath__49_0_I1817 (.Y(N6852), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[12]));
NOR2BX1 inst_cellmath__49_0_I1818 (.Y(N6798), .AN(inst_cellmath__45[14]), .B(inst_cellmath__45[15]));
XNOR2X1 inst_cellmath__50_0_I11060 (.Y(inst_cellmath__45[17]), .A(N6315), .B(N6188));
INVXL inst_cellmath__49_0_I1819 (.Y(N6819), .A(inst_cellmath__45[17]));
OAI21XL inst_cellmath__49_0_I1820 (.Y(N6840), .A0(inst_cellmath__45[16]), .A1(N6798), .B0(N6819));
NOR2X2 inst_cellmath__49_0_I1821 (.Y(N6765), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[14]));
NOR2X2 inst_cellmath__49_0_I1822 (.Y(N6787), .A(inst_cellmath__45[17]), .B(inst_cellmath__45[16]));
NOR2BX1 inst_cellmath__49_0_I1823 (.Y(N6827), .AN(inst_cellmath__45[18]), .B(inst_cellmath__45[19]));
INVXL inst_cellmath__49_0_I1824 (.Y(N6849), .A(inst_cellmath__45[21]));
OAI21XL inst_cellmath__49_0_I1825 (.Y(N6775), .A0(inst_cellmath__45[20]), .A1(N6827), .B0(N6849));
NOR2BXL inst_cellmath__49_0_I4579 (.Y(N6760), .AN(inst_cellmath__45[22]), .B(inst_cellmath__45[23]));
NOR2XL inst_cellmath__49_0_I4783 (.Y(N10869), .A(inst_cellmath__45[24]), .B(N6760));
OR2XL inst_cellmath__49_0_I11289 (.Y(N6804), .A(inst_cellmath__45[25]), .B(N10869));
NAND2BXL inst_cellmath__49_0_I1833 (.Y(N6842), .AN(N6774), .B(N6794));
OAI2BB1X1 inst_cellmath__49_0_I11290 (.Y(N6834), .A0N(N6802), .A1N(N6842), .B0(N6821));
NAND2X2 inst_cellmath__49_0_I1836 (.Y(N6810), .A(N6774), .B(N6794));
NAND2X2 inst_cellmath__49_0_I1837 (.Y(N6829), .A(N6802), .B(N6821));
NAND2BXL inst_cellmath__49_0_I1838 (.Y(N6777), .AN(N6832), .B(N6852));
INVXL inst_cellmath__49_0_I1839 (.Y(N6797), .A(N6787));
AOI21XL inst_cellmath__49_0_I1840 (.Y(N6818), .A0(N6765), .A1(N6777), .B0(N6797));
NAND2X4 inst_cellmath__49_0_I1841 (.Y(N6838), .A(N6832), .B(N6852));
NAND2X4 inst_cellmath__49_0_I1842 (.Y(N6762), .A(N6787), .B(N6765));
NAND2BXL inst_cellmath__49_0_I1843 (.Y(N6806), .AN(N6795), .B(N6816));
INVXL inst_cellmath__49_0_I1844 (.Y(N6825), .A(N6845));
AOI21XL inst_cellmath__49_0_I1845 (.Y(N6847), .A0(N6823), .A1(N6806), .B0(N6825));
NAND2BXL inst_cellmath__49_0_I1848 (.Y(N6782), .AN(N6829), .B(N6810));
NOR2X4 inst_cellmath__49_0_I1849 (.Y(N6768), .A(N6810), .B(N6829));
NOR2BX1 inst_cellmath__49_0_I1850 (.Y(N6811), .AN(N6838), .B(N6762));
INVXL inst_cellmath__49_0_I1851 (.Y(N6831), .A(N6793));
OAI21X1 inst_cellmath__49_0_I1852 (.Y(N6851), .A0(N6773), .A1(N6811), .B0(N6831));
NOR2X4 inst_cellmath__49_0_I1853 (.Y(N6779), .A(N6838), .B(N6762));
NAND2BX4 inst_cellmath__49_0_I1855 (.Y(N6839), .AN(N6763), .B(N6768));
INVX3 inst_cellmath__49_0_I1856 (.Y(N6764), .A(N6830));
AOI21X4 inst_cellmath__49_0_I1857 (.Y(inst_cellmath__49[3]), .A0(N6839), .A1(N6779), .B0(N6764));
NAND2XL inst_cellmath__49_0_I1858 (.Y(N6808), .A(N6768), .B(N6763));
NAND2X2 inst_cellmath__49_0_I1859 (.Y(N6778), .A(N6830), .B(N6779));
AOI21XL inst_cellmath__49_0_I1864 (.Y(N6800), .A0(N6830), .A1(N6818), .B0(N6847));
OAI21X1 inst_cellmath__49_0_I1865 (.Y(inst_cellmath__49[1]), .A0(N6778), .A1(N6834), .B0(N6800));
NOR2BX1 inst_cellmath__49_0_I1866 (.Y(N6785), .AN(inst_cellmath__45[0]), .B(inst_cellmath__45[1]));
OAI21XL inst_cellmath__49_0_I1867 (.Y(N6772), .A0(N6829), .A1(N6848), .B0(N6783));
OAI21XL inst_cellmath__49_0_I1868 (.Y(N6815), .A0(N6762), .A1(N6812), .B0(N6840));
OAI21X1 inst_cellmath__49_0_I1869 (.Y(N6855), .A0(N6793), .A1(N6775), .B0(N6804));
AOI21XL inst_cellmath__49_0_I1870 (.Y(N6801), .A0(N6768), .A1(N6785), .B0(N6772));
AOI21X1 inst_cellmath__49_0_I1871 (.Y(N6843), .A0(N6830), .A1(N6815), .B0(N6855));
OAI21X1 inst_cellmath__49_0_I1872 (.Y(inst_cellmath__49[0]), .A0(N6778), .A1(N6801), .B0(N6843));
NOR2XL inst_cellmath__71_1_I11001 (.Y(inst_cellmath__49[5]), .A(N6808), .B(N6778));
OR2XL cmpoi_A_I11458 (.Y(N17966), .A(a_sign), .B(b_sign));
AOI22XL cmpoi_A_I11459 (.Y(N645), .A0(inst_cellmath__6), .A1(N17966), .B0(a_sign), .B1(b_sign));
NAND2XL inst_cellmath__66_0_I1882 (.Y(N6958), .A(inst_cellmath__11), .B(inst_cellmath__16));
NOR2XL inst_cellmath__66_0_I1884 (.Y(inst_cellmath__66), .A(N645), .B(N6958));
INVXL inst_cellmath__64__48__2WWMM_I1885 (.Y(N7017), .A(a_sign));
INVXL inst_cellmath__64__48__2WWMM_I1909 (.Y(N7034), .A(inst_cellmath__18));
NOR2BX1 inst_cellmath__64__48__2WWMM_I4581 (.Y(N7050), .AN(N7034), .B(b_sign));
NAND2XL inst_cellmath__64__48__2WWMM_I1912 (.Y(N7004), .A(b_man[0]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1913 (.Y(N7064), .A(b_man[1]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1915 (.Y(N6987), .A(b_man[2]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1916 (.Y(N7045), .A(b_man[3]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1917 (.Y(N6969), .A(b_man[4]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1918 (.Y(N7028), .A(b_man[5]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1920 (.Y(N7086), .A(b_man[6]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1921 (.Y(N7011), .A(b_man[7]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1922 (.Y(N7071), .A(b_man[8]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1923 (.Y(N6995), .A(b_man[9]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1925 (.Y(N7054), .A(b_man[10]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1926 (.Y(N6977), .A(b_man[11]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1927 (.Y(N7035), .A(b_man[12]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1928 (.Y(N7092), .A(b_man[13]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1930 (.Y(N7016), .A(b_man[14]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1931 (.Y(N7076), .A(b_man[15]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1932 (.Y(N7000), .A(b_man[16]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1933 (.Y(N7060), .A(b_man[17]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1935 (.Y(N6984), .A(b_man[18]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1936 (.Y(N7042), .A(b_man[19]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1937 (.Y(N6966), .A(b_man[20]), .B(N7034));
NAND2XL inst_cellmath__64__48__2WWMM_I1938 (.Y(N7025), .A(b_man[21]), .B(N7034));
INVXL inst_cellmath__64__48__2WWMM_I1940 (.Y(N7090), .A(inst_cellmath__13));
INVXL inst_cellmath__64__48__2WWMM_I1941 (.Y(N7096), .A(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1943 (.Y(N710), .A0(N7050), .A1(N7096), .B0(N7017), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1944 (.Y(inst_cellmath__64[0]), .A0(N7096), .A1(N7004), .B0(N5224), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1945 (.Y(inst_cellmath__64[1]), .A0(N7064), .A1(N7096), .B0(N4820), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1946 (.Y(inst_cellmath__64[2]), .A0(N7096), .A1(N6987), .B0(N4338), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1947 (.Y(inst_cellmath__64[3]), .A0(N7096), .A1(N7045), .B0(N4801), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1948 (.Y(inst_cellmath__64[4]), .A0(N7096), .A1(N6969), .B0(N4866), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1949 (.Y(inst_cellmath__64[5]), .A0(N7096), .A1(N7028), .B0(N4934), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1950 (.Y(inst_cellmath__64[6]), .A0(N7096), .A1(N7086), .B0(N4847), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1952 (.Y(inst_cellmath__64[7]), .A0(N7096), .A1(N7011), .B0(N4912), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1953 (.Y(inst_cellmath__64[8]), .A0(N7096), .A1(N7071), .B0(N4829), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1954 (.Y(inst_cellmath__64[9]), .A0(N7096), .A1(N6995), .B0(N4893), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1955 (.Y(inst_cellmath__64[10]), .A0(N7096), .A1(N7054), .B0(N4807), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1956 (.Y(inst_cellmath__64[11]), .A0(N7096), .A1(N6977), .B0(N4875), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1957 (.Y(inst_cellmath__64[12]), .A0(N7096), .A1(N7035), .B0(N4791), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1958 (.Y(inst_cellmath__64[13]), .A0(N7096), .A1(N7092), .B0(N4854), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1959 (.Y(inst_cellmath__64[14]), .A0(N7096), .A1(N7016), .B0(N4922), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1961 (.Y(inst_cellmath__64[15]), .A0(N7096), .A1(N7076), .B0(N4839), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1962 (.Y(inst_cellmath__64[16]), .A0(N7096), .A1(N7000), .B0(N4901), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1963 (.Y(inst_cellmath__64[17]), .A0(N7096), .A1(N7060), .B0(N4817), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1964 (.Y(inst_cellmath__64[18]), .A0(N7096), .A1(N6984), .B0(N4884), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1965 (.Y(inst_cellmath__64[19]), .A0(N7096), .A1(N7042), .B0(N4796), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1966 (.Y(inst_cellmath__64[20]), .A0(N7096), .A1(N6966), .B0(N4864), .B1(N7090));
AOI22XL inst_cellmath__64__48__2WWMM_I1967 (.Y(inst_cellmath__64[21]), .A0(N7096), .A1(N7025), .B0(N4931), .B1(N7090));
MXI2XL inst_cellmath__67_0_I1968 (.Y(N7182), .A(inst_cellmath__66), .B(N710), .S0(inst_cellmath__63));
NOR2XL inst_cellmath__67_0_I1969 (.Y(N7191), .A(inst_cellmath__63), .B(N706));
MXI2XL inst_cellmath__67_0_I11293 (.Y(N7185), .A(inst_cellmath__48), .B(inst_cellmath__6), .S0(inst_cellmath__49[5]));
MXI2XL inst_cellmath__67_0_I1971 (.Y(x[31]), .A(N7182), .B(N7185), .S0(N7191));
CLKINVX4 inst_cellmath__50_0_I1972 (.Y(N7197), .A(inst_cellmath__49[3]));
CLKINVX8 inst_cellmath__50_0_I4428 (.Y(N10733), .A(N7197));
NOR2BX2 inst_cellmath__50_0_I11061 (.Y(N17663), .AN(N6808), .B(N6778));
OAI21X2 inst_cellmath__50_0_I11062 (.Y(N17620), .A0(N6778), .A1(N6782), .B0(N6851));
INVXL inst_cellmath__50_0_I11063 (.Y(N17653), .A(N10733));
CLKAND2X3 inst_cellmath__50_0_I11064 (.Y(N7284), .A(inst_cellmath__45[1]), .B(N17653));
INVX2 inst_cellmath__50_0_I11065 (.Y(N10736), .A(N10733));
NAND2BXL inst_cellmath__50_0_I11297 (.Y(N17618), .AN(N10736), .B(inst_cellmath__45[5]));
NAND2XL inst_cellmath__50_0_I11070 (.Y(N17664), .A(N10736), .B(inst_cellmath__45[13]));
MX2XL inst_cellmath__50_0_I11298 (.Y(N17644), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[13]), .S0(N10736));
INVX3 inst_cellmath__50_0_I11072 (.Y(N10737), .A(N10733));
INVXL inst_cellmath__50_0_I11074 (.Y(N17660), .A(inst_cellmath__45[9]));
OR2XL inst_cellmath__50_0_I11374 (.Y(N17638), .A(N17660), .B(N10737));
NAND2XL inst_cellmath__50_0_I11077 (.Y(N17628), .A(N10737), .B(inst_cellmath__45[17]));
MX2XL inst_cellmath__50_0_I11302 (.Y(N17655), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[17]), .S0(N10737));
CLKINVX8 inst_cellmath__50_0_I11079 (.Y(N7234), .A(N17663));
AOI21XL inst_cellmath__50_0_I11080 (.Y(N17642), .A0(N17664), .A1(N17618), .B0(N17663));
NAND2X1 inst_cellmath__50_0_I11081 (.Y(N7319), .A(N7234), .B(N17644));
AOI21XL inst_cellmath__50_0_I11082 (.Y(N17632), .A0(N17628), .A1(N17638), .B0(N17663));
NAND2XL inst_cellmath__50_0_I11083 (.Y(N17626), .A(inst_cellmath__45[1]), .B(N17653));
NOR2XL inst_cellmath__50_0_I11084 (.Y(N17649), .A(N7234), .B(N17626));
MXI2XL inst_cellmath__50_0_I11085 (.Y(N7240), .A(N7284), .B(N17655), .S0(N7234));
INVX3 inst_cellmath__50_0_I11086 (.Y(N17637), .A(N17620));
CLKINVX12 inst_cellmath__50_0_I11087 (.Y(N7286), .A(N17637));
INVXL buf1_A_I11460 (.Y(N17974), .A(N17637));
INVXL buf1_A_I11461 (.Y(N7272), .A(N17974));
NOR2XL inst_cellmath__50_0_I11089 (.Y(N17631), .A(N17642), .B(N7272));
NOR3XL inst_cellmath__50_0_I11303 (.Y(N17648), .A(N17620), .B(N17632), .C(N17649));
NOR2X1 inst_cellmath__50_0_I11092 (.Y(N7253), .A(N17631), .B(N17648));
INVX2 inst_cellmath__50_0_I4433 (.Y(N10738), .A(N10733));
INVX2 inst_cellmath__50_0_I4430 (.Y(N10735), .A(N10733));
INVX2 inst_cellmath__50_0_I4429 (.Y(N10734), .A(N10733));
CLKAND2X2 inst_cellmath__50_0_I1973 (.Y(N7211), .A(N7197), .B(inst_cellmath__45[0]));
CLKAND2X3 inst_cellmath__50_0_I1975 (.Y(N7357), .A(inst_cellmath__45[2]), .B(N10738));
AND2XL inst_cellmath__50_0_I1976 (.Y(N7263), .A(inst_cellmath__45[3]), .B(N10734));
AND2XL inst_cellmath__50_0_I1977 (.Y(N7335), .A(inst_cellmath__45[4]), .B(N10734));
AND2XL inst_cellmath__50_0_I1978 (.Y(N7242), .A(N10735), .B(inst_cellmath__45[5]));
AND2XL inst_cellmath__50_0_I1979 (.Y(N7316), .A(N10735), .B(inst_cellmath__45[6]));
AND2XL inst_cellmath__50_0_I1980 (.Y(N7221), .A(N10735), .B(inst_cellmath__45[7]));
MX2XL inst_cellmath__50_0_I1981 (.Y(N7294), .A(inst_cellmath__45[0]), .B(inst_cellmath__45[8]), .S0(N10735));
MX2XL inst_cellmath__50_0_I1982 (.Y(N7331), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[9]), .S0(N10735));
MX2XL inst_cellmath__50_0_I1983 (.Y(N7199), .A(inst_cellmath__45[2]), .B(inst_cellmath__45[10]), .S0(N10736));
MX2XL inst_cellmath__50_0_I1984 (.Y(N7236), .A(inst_cellmath__45[3]), .B(inst_cellmath__45[11]), .S0(N10736));
MX2XL inst_cellmath__50_0_I1985 (.Y(N7273), .A(inst_cellmath__45[4]), .B(inst_cellmath__45[12]), .S0(N10736));
MX2XL inst_cellmath__50_0_I1987 (.Y(N7345), .A(inst_cellmath__45[6]), .B(inst_cellmath__45[14]), .S0(N10736));
MX2XL inst_cellmath__50_0_I1988 (.Y(N7216), .A(inst_cellmath__45[7]), .B(inst_cellmath__45[15]), .S0(N10737));
OR2XL inst_cellmath__50_0_I4698 (.Y(N10721), .A(inst_cellmath__45[8]), .B(N10734));
NAND2BX1 inst_cellmath__50_0_I4699 (.Y(N10715), .AN(inst_cellmath__45[16]), .B(N10734));
CLKAND2X2 inst_cellmath__50_0_I4454 (.Y(N7252), .A(N10715), .B(N10721));
MX2XL inst_cellmath__50_0_I1991 (.Y(N7323), .A(inst_cellmath__45[10]), .B(inst_cellmath__45[18]), .S0(N10737));
MX2XL inst_cellmath__50_0_I1992 (.Y(N7360), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[19]), .S0(N10737));
MX2XL inst_cellmath__50_0_I1993 (.Y(N7229), .A(inst_cellmath__45[12]), .B(inst_cellmath__45[20]), .S0(N10737));
MX2XL inst_cellmath__50_0_I1994 (.Y(N7267), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[21]), .S0(N10738));
MX2XL inst_cellmath__50_0_I1995 (.Y(N7304), .A(inst_cellmath__45[14]), .B(inst_cellmath__45[22]), .S0(N10738));
MX2XL inst_cellmath__50_0_I1996 (.Y(N7340), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[23]), .S0(N10738));
MX2XL inst_cellmath__50_0_I1997 (.Y(N7208), .A(inst_cellmath__45[16]), .B(inst_cellmath__45[24]), .S0(N10738));
NAND2X4 inst_cellmath__50_0_I1999 (.Y(N7204), .A(N7234), .B(N7211));
NAND2X4 inst_cellmath__50_0_I2000 (.Y(N7279), .A(N7234), .B(N7284));
NAND2X2 inst_cellmath__50_0_I2001 (.Y(N7351), .A(N7234), .B(N7357));
NAND2XL inst_cellmath__50_0_I2002 (.Y(N7257), .A(N7263), .B(N7234));
NAND2XL inst_cellmath__50_0_I2003 (.Y(N7329), .A(N7335), .B(N7234));
NAND2XL inst_cellmath__50_0_I2004 (.Y(N7235), .A(N7242), .B(N7234));
NAND2XL inst_cellmath__50_0_I2005 (.Y(N7308), .A(N7316), .B(N7234));
NAND2XL inst_cellmath__50_0_I2006 (.Y(N7214), .A(N7221), .B(N7234));
NAND2X1 inst_cellmath__50_0_I2007 (.Y(N7287), .A(N7234), .B(N7294));
NAND2X1 inst_cellmath__50_0_I2008 (.Y(N7359), .A(N7234), .B(N7331));
NAND2X1 inst_cellmath__50_0_I2009 (.Y(N7265), .A(N7234), .B(N7199));
NAND2X1 inst_cellmath__50_0_I2010 (.Y(N7339), .A(N7234), .B(N7236));
NAND2X1 inst_cellmath__50_0_I2011 (.Y(N7246), .A(N7234), .B(N7273));
NAND2X1 inst_cellmath__50_0_I2013 (.Y(N7225), .A(N7234), .B(N7345));
NAND2X1 inst_cellmath__50_0_I2014 (.Y(N7298), .A(N7234), .B(N7216));
MXI2X1 inst_cellmath__50_0_I2015 (.Y(N7202), .A(N7211), .B(N7252), .S0(N7234));
MXI2X1 inst_cellmath__50_0_I2017 (.Y(N7277), .A(N7357), .B(N7323), .S0(N7234));
MXI2X1 inst_cellmath__50_0_I2018 (.Y(N7313), .A(N7263), .B(N7360), .S0(N7234));
MXI2X1 inst_cellmath__50_0_I2019 (.Y(N7349), .A(N7335), .B(N7229), .S0(N7234));
MXI2XL inst_cellmath__50_0_I2020 (.Y(N7219), .A(N7242), .B(N7267), .S0(N7234));
MXI2XL inst_cellmath__50_0_I2021 (.Y(N7255), .A(N7316), .B(N7304), .S0(N7234));
MXI2XL inst_cellmath__50_0_I2022 (.Y(N7292), .A(N7221), .B(N7340), .S0(N7234));
MXI2XL inst_cellmath__50_0_I2023 (.Y(N7327), .A(N7294), .B(N7208), .S0(N7234));
NOR2X4 inst_cellmath__50_0_I2028 (.Y(N7322), .A(N7286), .B(N7204));
NOR2X2 inst_cellmath__50_0_I2029 (.Y(N7228), .A(N7286), .B(N7279));
NOR2X2 inst_cellmath__50_0_I2030 (.Y(N7301), .A(N7286), .B(N7351));
NOR2XL inst_cellmath__50_0_I2031 (.Y(N7207), .A(N7257), .B(N7286));
MXI2XL inst_cellmath__50_0_I2032 (.Y(N7282), .A(N7329), .B(N7204), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2033 (.Y(N7317), .A(N7235), .B(N7279), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2034 (.Y(N7354), .A(N7308), .B(N7351), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2035 (.Y(N7224), .A(N7214), .B(N7257), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2036 (.Y(N7261), .A(N7287), .B(N7329), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2037 (.Y(N7297), .A(N7359), .B(N7235), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2038 (.Y(N7333), .A(N7265), .B(N7308), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2039 (.Y(N7200), .A(N7339), .B(N7214), .S0(N7286));
MXI2X1 inst_cellmath__50_0_I2040 (.Y(N7238), .A(N7246), .B(N7287), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2041 (.Y(N7276), .A(N7319), .B(N7359), .S0(N7286));
MXI2X1 inst_cellmath__50_0_I2042 (.Y(N7312), .A(N7225), .B(N7265), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2043 (.Y(N7348), .A(N7298), .B(N7339), .S0(N7286));
MXI2X1 inst_cellmath__50_0_I2044 (.Y(N7218), .A(N7202), .B(N7246), .S0(N7286));
MXI2X1 inst_cellmath__50_0_I2046 (.Y(N7290), .A(N7277), .B(N7225), .S0(N7286));
MXI2X1 inst_cellmath__50_0_I2047 (.Y(N7326), .A(N7313), .B(N7298), .S0(N7286));
MXI2X1 inst_cellmath__50_0_I2048 (.Y(N7363), .A(N7349), .B(N7202), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2049 (.Y(N7232), .A(N7219), .B(N7240), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2050 (.Y(N7269), .A(N7255), .B(N7277), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2051 (.Y(N7305), .A(N7292), .B(N7313), .S0(N7286));
MXI2XL inst_cellmath__50_0_I2052 (.Y(N7342), .A(N7327), .B(N7349), .S0(N7286));
CLKINVX6 inst_cellmath__50_0_I2053 (.Y(N7206), .A(inst_cellmath__49[0]));
NAND2X4 inst_cellmath__50_0_I2056 (.Y(N7336), .A(N7322), .B(N7206));
MXI2XL inst_cellmath__50_0_I2057 (.Y(N7244), .A(N7322), .B(N7228), .S0(N7206));
MXI2X1 inst_cellmath__50_0_I2058 (.Y(N7280), .A(N7228), .B(N7301), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2059 (.Y(N7315), .A(N7301), .B(N7207), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2060 (.Y(N7352), .A(N7207), .B(N7282), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2061 (.Y(N7222), .A(N7282), .B(N7317), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2062 (.Y(N7258), .A(N7317), .B(N7354), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2063 (.Y(N7295), .A(N7354), .B(N7224), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2064 (.Y(N7330), .A(N7224), .B(N7261), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2065 (.Y(N7198), .A(N7261), .B(N7297), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2066 (.Y(N7237), .A(N7297), .B(N7333), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2067 (.Y(N7274), .A(N7333), .B(N7200), .S0(N7206));
MXI2X1 inst_cellmath__50_0_I2068 (.Y(N7310), .A(N7200), .B(N7238), .S0(N7206));
MXI2X1 inst_cellmath__50_0_I2069 (.Y(N7346), .A(N7238), .B(N7276), .S0(N7206));
MXI2X1 inst_cellmath__50_0_I2070 (.Y(N7215), .A(N7276), .B(N7312), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2071 (.Y(N7251), .A(N7312), .B(N7348), .S0(N7206));
MXI2X1 inst_cellmath__50_0_I2072 (.Y(N7289), .A(N7348), .B(N7218), .S0(N7206));
MXI2X1 inst_cellmath__50_0_I2073 (.Y(N7324), .A(N7218), .B(N7253), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2074 (.Y(N7361), .A(N7253), .B(N7290), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2075 (.Y(N7230), .A(N7290), .B(N7326), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2076 (.Y(N7266), .A(N7326), .B(N7363), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2077 (.Y(N7303), .A(N7363), .B(N7232), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2078 (.Y(N7341), .A(N7232), .B(N7269), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2079 (.Y(N7209), .A(N7269), .B(N7305), .S0(N7206));
MXI2XL inst_cellmath__50_0_I2080 (.Y(N7247), .A(N7305), .B(N7342), .S0(N7206));
INVX2 inst_cellmath__50_0_I2081 (.Y(N7243), .A(inst_cellmath__49[1]));
CLKINVX4 inst_cellmath__50_0_I2082 (.Y(N7260), .A(N7243));
NOR2XL inst_cellmath__50_0_I2085 (.Y(inst_cellmath__50[1]), .A(N7260), .B(N7244));
MXI2X1 inst_cellmath__50_0_I2086 (.Y(inst_cellmath__50[2]), .A(N7280), .B(N7336), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2087 (.Y(inst_cellmath__50[3]), .A(N7315), .B(N7244), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2088 (.Y(inst_cellmath__50[4]), .A(N7352), .B(N7280), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2089 (.Y(inst_cellmath__50[5]), .A(N7222), .B(N7315), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2090 (.Y(inst_cellmath__50[6]), .A(N7258), .B(N7352), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2091 (.Y(inst_cellmath__50[7]), .A(N7295), .B(N7222), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2092 (.Y(inst_cellmath__50[8]), .A(N7330), .B(N7258), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2093 (.Y(inst_cellmath__50[9]), .A(N7198), .B(N7295), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2094 (.Y(inst_cellmath__50[10]), .A(N7237), .B(N7330), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2095 (.Y(inst_cellmath__50[11]), .A(N7274), .B(N7198), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2096 (.Y(inst_cellmath__50[12]), .A(N7310), .B(N7237), .S0(N7260));
MXI2X1 inst_cellmath__50_0_I2097 (.Y(inst_cellmath__50[13]), .A(N7346), .B(N7274), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2098 (.Y(inst_cellmath__50[14]), .A(N7215), .B(N7310), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2099 (.Y(inst_cellmath__50[15]), .A(N7251), .B(N7346), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2100 (.Y(inst_cellmath__50[16]), .A(N7289), .B(N7215), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2101 (.Y(inst_cellmath__50[17]), .A(N7324), .B(N7251), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2102 (.Y(inst_cellmath__50[18]), .A(N7361), .B(N7289), .S0(N7260));
MXI2X1 inst_cellmath__50_0_I2103 (.Y(inst_cellmath__50[19]), .A(N7230), .B(N7324), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2104 (.Y(inst_cellmath__50[20]), .A(N7266), .B(N7361), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2105 (.Y(inst_cellmath__50[21]), .A(N7303), .B(N7230), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2106 (.Y(inst_cellmath__50[22]), .A(N7341), .B(N7266), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2107 (.Y(inst_cellmath__50[23]), .A(N7209), .B(N7303), .S0(N7260));
MXI2XL inst_cellmath__50_0_I2108 (.Y(inst_cellmath__50[24]), .A(N7247), .B(N7341), .S0(N7260));
INVXL buf1_A_I4745 (.Y(N10790), .A(inst_cellmath__50[2]));
INVXL buf1_A_I4746 (.Y(N2855), .A(N10790));
INVXL inst_cellmath__43__26__I2109 (.Y(N7503), .A(inst_cellmath__33[24]));
XNOR2X1 inst_cellmath__43__26__I4589 (.Y(N626), .A(N7503), .B(N1693));
NAND2BXL cynw_cm_float_add2_ieee_I4590 (.Y(N627), .AN(inst_cellmath__30), .B(N626));
OAI21XL cynw_cm_float_add2_ieee_I4591 (.Y(N7524), .A0(inst_cellmath__33[24]), .A1(N1693), .B0(inst_cellmath__30));
AND2XL cynw_cm_float_add2_ieee_I2119 (.Y(N7530), .A(N7524), .B(N627));
AOI22XL cynw_cm_float_add2_ieee_I2124 (.Y(inst_cellmath__43), .A0(N5967), .A1(N7503), .B0(N7530), .B1(inst_cellmath__39[25]));
MX2XL cynw_cm_float_add2_ieee_I2127 (.Y(inst_cellmath__53), .A(inst_cellmath__50[1]), .B(inst_cellmath__43), .S0(inst_cellmath__49[1]));
INVXL inst_cellmath__5_0_I2128 (.Y(N7558), .A(rm[1]));
AND3XL inst_cellmath__5_0_I4592 (.Y(inst_cellmath__5), .A(rm[0]), .B(N4582), .C(N7558));
INVXL inst_cellmath__55__39__I2132 (.Y(N7567), .A(inst_cellmath__5));
NOR2XL inst_cellmath__55__39__I2133 (.Y(N635), .A(N7567), .B(inst_cellmath__48));
AND2XL cynw_cm_float_add2_ieee_I2134 (.Y(N634), .A(inst_cellmath__6), .B(inst_cellmath__48));
AND3XL cynw_cm_float_add2_ieee_I4593 (.Y(inst_cellmath__8), .A(rm[2]), .B(N7558), .C(N4581));
AND3XL cynw_cm_float_add2_ieee_I4594 (.Y(inst_cellmath__4), .A(N4581), .B(N4582), .C(N7558));
NOR2XL inst_cellmath__54__33__I2144 (.Y(N7603), .A(inst_cellmath__43), .B(N1693));
OAI21X2 inst_cellmath__54__33__I4398 (.Y(N7606), .A0(N7260), .A1(N7336), .B0(N7603));
MX2XL cynw_cm_float_add2_ieee_I2149 (.Y(inst_cellmath__54), .A(N7606), .B(N1693), .S0(inst_cellmath__49[1]));
OAI21X1 cynw_cm_float_add2_ieee_I4399 (.Y(N7625), .A0(inst_cellmath__50[2]), .A1(inst_cellmath__54), .B0(inst_cellmath__4));
NOR3XL cynw_cm_float_add2_ieee_I4595 (.Y(N7640), .A(inst_cellmath__8), .B(N635), .C(N634));
OAI2BB1XL cynw_cm_float_add2_ieee_I4473 (.Y(N7647), .A0N(N7640), .A1N(N7625), .B0(inst_cellmath__53));
OAI21XL cynw_cm_float_add2_ieee_I4704 (.Y(N639), .A0(N635), .A1(N634), .B0(inst_cellmath__54));
AND2X1 inst_cellmath__55_0_I2164 (.Y(N7661), .A(N7647), .B(N639));
INVX2 inst_cellmath__55_0_I2165 (.Y(inst_cellmath__55), .A(N7661));
CLKAND2X6 inst_cellmath__57_0_I2168 (.Y(N7732), .A(N2855), .B(inst_cellmath__55));
AND2XL inst_cellmath__57_0_I2169 (.Y(N7708), .A(inst_cellmath__50[3]), .B(inst_cellmath__55));
AND2X2 inst_cellmath__57_0_I2170 (.Y(N7772), .A(inst_cellmath__50[4]), .B(inst_cellmath__50[3]));
AND2XL inst_cellmath__57_0_I2171 (.Y(N7693), .A(inst_cellmath__50[5]), .B(inst_cellmath__50[4]));
AND2X1 inst_cellmath__57_0_I2172 (.Y(N7757), .A(inst_cellmath__50[5]), .B(inst_cellmath__50[6]));
AND2XL inst_cellmath__57_0_I2173 (.Y(N7671), .A(inst_cellmath__50[7]), .B(inst_cellmath__50[6]));
AND2X1 inst_cellmath__57_0_I2174 (.Y(N7741), .A(inst_cellmath__50[8]), .B(inst_cellmath__50[7]));
AND2XL inst_cellmath__57_0_I2175 (.Y(N7796), .A(inst_cellmath__50[8]), .B(inst_cellmath__50[9]));
CLKAND2X2 inst_cellmath__57_0_I2176 (.Y(N7718), .A(inst_cellmath__50[10]), .B(inst_cellmath__50[9]));
AND2XL inst_cellmath__57_0_I2177 (.Y(N7782), .A(inst_cellmath__50[11]), .B(inst_cellmath__50[10]));
CLKAND2X2 inst_cellmath__57_0_I2178 (.Y(N7702), .A(inst_cellmath__50[12]), .B(inst_cellmath__50[11]));
AND2XL inst_cellmath__57_0_I2179 (.Y(N7763), .A(inst_cellmath__50[12]), .B(inst_cellmath__50[13]));
CLKAND2X2 inst_cellmath__57_0_I2180 (.Y(N7682), .A(inst_cellmath__50[14]), .B(inst_cellmath__50[13]));
AND2XL inst_cellmath__57_0_I2181 (.Y(N7747), .A(inst_cellmath__50[15]), .B(inst_cellmath__50[14]));
CLKAND2X2 inst_cellmath__57_0_I2182 (.Y(N7801), .A(inst_cellmath__50[16]), .B(inst_cellmath__50[15]));
AND2XL inst_cellmath__57_0_I2183 (.Y(N7728), .A(inst_cellmath__50[16]), .B(inst_cellmath__50[17]));
CLKAND2X2 inst_cellmath__57_0_I2184 (.Y(N7788), .A(inst_cellmath__50[18]), .B(inst_cellmath__50[17]));
AND2XL inst_cellmath__57_0_I2185 (.Y(N7705), .A(inst_cellmath__50[19]), .B(inst_cellmath__50[18]));
CLKAND2X2 inst_cellmath__57_0_I2186 (.Y(N7769), .A(inst_cellmath__50[19]), .B(inst_cellmath__50[20]));
AND2XL inst_cellmath__57_0_I2187 (.Y(N7688), .A(inst_cellmath__50[20]), .B(inst_cellmath__50[21]));
CLKAND2X2 inst_cellmath__57_0_I2188 (.Y(N7754), .A(inst_cellmath__50[21]), .B(inst_cellmath__50[22]));
CLKAND2X2 inst_cellmath__57_0_I2189 (.Y(N7737), .A(inst_cellmath__50[23]), .B(inst_cellmath__50[24]));
INVXL inst_cellmath__57_0_I2190 (.Y(N7712), .A(N2855));
INVXL inst_cellmath__57_0_I2191 (.Y(N7748), .A(N7732));
NAND2XL inst_cellmath__57_0_I2192 (.Y(N7751), .A(N7708), .B(N2855));
NAND2X8 inst_cellmath__57_0_I2193 (.Y(N7699), .A(N7772), .B(N7732));
NAND2XL inst_cellmath__57_0_I2194 (.Y(N7678), .A(N7693), .B(N7708));
NAND2XL inst_cellmath__57_0_I2195 (.Y(N7746), .A(N7757), .B(N7772));
NAND2XL inst_cellmath__57_0_I2196 (.Y(N7800), .A(N7671), .B(N7693));
NAND2X4 inst_cellmath__57_0_I2197 (.Y(N7724), .A(N7757), .B(N7741));
NAND2XL inst_cellmath__57_0_I2198 (.Y(N7786), .A(N7796), .B(N7671));
NAND2XL inst_cellmath__57_0_I2199 (.Y(N7704), .A(N7718), .B(N7741));
NAND2XL inst_cellmath__57_0_I2200 (.Y(N7766), .A(N7782), .B(N7796));
NAND2X4 inst_cellmath__57_0_I2201 (.Y(N7686), .A(N7718), .B(N7702));
NAND2XL inst_cellmath__57_0_I2202 (.Y(N7753), .A(N7763), .B(N7782));
NAND2XL inst_cellmath__57_0_I2203 (.Y(N7808), .A(N7682), .B(N7702));
NAND2XL inst_cellmath__57_0_I2204 (.Y(N7735), .A(N7747), .B(N7763));
NAND2X4 inst_cellmath__57_0_I2205 (.Y(N7792), .A(N7682), .B(N7801));
NAND2XL inst_cellmath__57_0_I2206 (.Y(N7710), .A(N7728), .B(N7747));
NAND2XL inst_cellmath__57_0_I2207 (.Y(N7775), .A(N7801), .B(N7788));
NAND2XL inst_cellmath__57_0_I2208 (.Y(N7695), .A(N7705), .B(N7728));
NAND2X4 inst_cellmath__57_0_I2209 (.Y(N7759), .A(N7769), .B(N7788));
NAND3XL inst_cellmath__57_0_I2212 (.Y(N7798), .A(N7688), .B(inst_cellmath__50[22]), .C(inst_cellmath__50[23]));
NAND2X4 inst_cellmath__57_0_I2213 (.Y(N7721), .A(N7737), .B(N7754));
INVXL inst_cellmath__57_0_I2214 (.Y(N7776), .A(N7712));
INVXL inst_cellmath__57_0_I2215 (.Y(N7803), .A(N7748));
INVXL inst_cellmath__57_0_I2216 (.Y(N7696), .A(N7751));
INVXL inst_cellmath__57_0_I2217 (.Y(N7729), .A(N7699));
NOR2XL inst_cellmath__57_0_I2218 (.Y(N7713), .A(N7678), .B(N7712));
NOR2XL inst_cellmath__57_0_I2219 (.Y(N7804), .A(N7746), .B(N7748));
NOR2XL inst_cellmath__57_0_I2220 (.Y(N7761), .A(N7800), .B(N7751));
NOR2X6 inst_cellmath__57_0_I2221 (.Y(N7706), .A(N7724), .B(N7699));
NOR2XL inst_cellmath__57_0_I2222 (.Y(N7691), .A(N7786), .B(N7678));
NOR2XL inst_cellmath__57_0_I2223 (.Y(N7755), .A(N7704), .B(N7746));
NOR2XL inst_cellmath__57_0_I2224 (.Y(N7668), .A(N7766), .B(N7800));
NOR2XL inst_cellmath__57_0_I2225 (.Y(N7739), .A(N7686), .B(N7724));
NOR2XL inst_cellmath__57_0_I2226 (.Y(N7795), .A(N7753), .B(N7786));
NOR2XL inst_cellmath__57_0_I2227 (.Y(N7717), .A(N7808), .B(N7704));
NOR2XL inst_cellmath__57_0_I2228 (.Y(N7781), .A(N7735), .B(N7766));
NOR2X4 inst_cellmath__57_0_I2229 (.Y(N7701), .A(N7792), .B(N7686));
NAND4BXL inst_cellmath__57_0_I11311 (.Y(N7758), .AN(N7710), .B(N7688), .C(N7795), .D(N7705));
NAND4BXL inst_cellmath__57_0_I11312 (.Y(N7672), .AN(N7775), .B(N7769), .C(N7717), .D(N7754));
NOR2X4 inst_cellmath__57_0_I2233 (.Y(N7768), .A(N7759), .B(N7721));
INVXL inst_cellmath__57_0_I2234 (.Y(N7676), .A(N7803));
INVXL inst_cellmath__57_0_I2235 (.Y(N7689), .A(N7713));
INVXL inst_cellmath__57_0_I2236 (.Y(N7722), .A(N7804));
INVX4 inst_cellmath__57_0_I2237 (.Y(N7667), .A(N7706));
NAND2XL inst_cellmath__57_0_I2238 (.Y(N7675), .A(N7755), .B(N7803));
NAND2XL inst_cellmath__57_0_I2239 (.Y(N7716), .A(N7781), .B(N7761));
NAND2XL inst_cellmath__57_0_I2240 (.Y(N7806), .A(N7701), .B(N7706));
NOR3BXL inst_cellmath__57_0_I2241 (.Y(N7791), .AN(N7691), .B(N7710), .C(N7753));
NOR4BX1 node_cs_const1_cs_A_I11314 (.Y(N10829), .AN(N7755), .B(N7775), .C(N7676), .D(N7808));
NOR3BXL inst_cellmath__57_0_I2243 (.Y(N7773), .AN(N7668), .B(N7695), .C(N7735));
NOR3BXL inst_cellmath__57_0_I2244 (.Y(N7694), .AN(N7739), .B(N7792), .C(N7759));
NOR3BXL inst_cellmath__57_0_I2247 (.Y(N7742), .AN(N7781), .B(N7695), .C(N7798));
NAND2X4 inst_cellmath__57_0_I2248 (.Y(N7797), .A(N7701), .B(N7768));
NAND2XL inst_cellmath__57_0_I2254 (.Y(N7684), .A(N7791), .B(N7776));
NAND2XL inst_cellmath__57_0_I2256 (.Y(N7731), .A(N7773), .B(N7696));
NAND2XL inst_cellmath__57_0_I2257 (.Y(N7679), .A(N7694), .B(N7729));
NAND2XL inst_cellmath__57_0_I2260 (.Y(N7670), .A(N7742), .B(N7761));
XNOR2X1 inst_cellmath__57_0_I2262 (.Y(inst_cellmath__57[0]), .A(inst_cellmath__55), .B(N7776));
XNOR2X1 inst_cellmath__57_0_I2263 (.Y(inst_cellmath__57[1]), .A(inst_cellmath__50[3]), .B(N7676));
XNOR2X1 inst_cellmath__57_0_I2264 (.Y(inst_cellmath__57[2]), .A(N7696), .B(inst_cellmath__50[4]));
XNOR2X1 inst_cellmath__57_0_I2265 (.Y(inst_cellmath__57[3]), .A(N7729), .B(inst_cellmath__50[5]));
XNOR2X1 inst_cellmath__57_0_I2266 (.Y(inst_cellmath__57[4]), .A(inst_cellmath__50[6]), .B(N7689));
XNOR2X1 inst_cellmath__57_0_I2267 (.Y(inst_cellmath__57[5]), .A(N7722), .B(inst_cellmath__50[7]));
XNOR2X1 inst_cellmath__57_0_I2268 (.Y(inst_cellmath__57[6]), .A(N7761), .B(inst_cellmath__50[8]));
XNOR2X1 inst_cellmath__57_0_I2269 (.Y(inst_cellmath__57[7]), .A(N7667), .B(inst_cellmath__50[9]));
NAND2XL node_cs_const1_cs_ii_A_I4747 (.Y(N10794), .A(N7691), .B(N7776));
XOR2XL node_cs_const1_cs_ii_A_I4748 (.Y(inst_cellmath__57[8]), .A(inst_cellmath__50[10]), .B(N10794));
XNOR2X1 inst_cellmath__57_0_I2271 (.Y(inst_cellmath__57[9]), .A(inst_cellmath__50[11]), .B(N7675));
NAND2XL node_cs_const1_cs_ii_A_I4749 (.Y(N10801), .A(N7668), .B(N7696));
XOR2XL node_cs_const1_cs_ii_A_I4750 (.Y(inst_cellmath__57[10]), .A(inst_cellmath__50[12]), .B(N10801));
NAND2XL node_cs_const1_cs_ii_A_I4751 (.Y(N10808), .A(N7739), .B(N7729));
XOR2XL node_cs_const1_cs_ii_A_I4752 (.Y(inst_cellmath__57[11]), .A(inst_cellmath__50[13]), .B(N10808));
NAND2XL node_cs_const1_cs_ii_A_I4753 (.Y(N10815), .A(N7795), .B(N7713));
XOR2XL node_cs_const1_cs_ii_A_I4754 (.Y(inst_cellmath__57[12]), .A(inst_cellmath__50[14]), .B(N10815));
NAND2XL node_cs_const1_cs_ii_A_I4755 (.Y(N10822), .A(N7717), .B(N7804));
XOR2XL node_cs_const1_cs_ii_A_I4756 (.Y(inst_cellmath__57[13]), .A(inst_cellmath__50[15]), .B(N10822));
XNOR2X1 inst_cellmath__57_0_I2276 (.Y(inst_cellmath__57[14]), .A(inst_cellmath__50[16]), .B(N7716));
XNOR2X1 inst_cellmath__57_0_I2277 (.Y(inst_cellmath__57[15]), .A(inst_cellmath__50[17]), .B(N7806));
XNOR2X1 inst_cellmath__57_0_I2278 (.Y(inst_cellmath__57[16]), .A(inst_cellmath__50[18]), .B(N7684));
XNOR2X1 node_cs_const1_cs_A_I4758 (.Y(inst_cellmath__57[17]), .A(inst_cellmath__50[19]), .B(N10829));
XNOR2X1 inst_cellmath__57_0_I2280 (.Y(inst_cellmath__57[18]), .A(inst_cellmath__50[20]), .B(N7731));
XNOR2X1 inst_cellmath__57_0_I2281 (.Y(inst_cellmath__57[19]), .A(inst_cellmath__50[21]), .B(N7679));
NOR2XL node_cs_const1_cs_A_I4759 (.Y(N10836), .A(N7758), .B(N7689));
XNOR2X1 node_cs_const1_cs_A_I4760 (.Y(inst_cellmath__57[20]), .A(inst_cellmath__50[22]), .B(N10836));
NOR2XL node_cs_const1_cs_A_I4761 (.Y(N10843), .A(N7672), .B(N7722));
XNOR2X1 node_cs_const1_cs_A_I4762 (.Y(inst_cellmath__57[21]), .A(inst_cellmath__50[23]), .B(N10843));
XNOR2X1 inst_cellmath__57_0_I2284 (.Y(inst_cellmath__57[22]), .A(N7670), .B(inst_cellmath__50[24]));
NOR2X4 inst_cellmath__59_0_I11214 (.Y(N17525), .A(N7797), .B(N7667));
INVXL buf1_A_I11462 (.Y(N17979), .A(N17525));
INVXL buf1_A_I11463 (.Y(inst_cellmath__57[23]), .A(N17979));
AOI21XL cynw_cm_float_add2_ieee_I11317 (.Y(N642), .A0(inst_cellmath__57[23]), .A1(inst_cellmath__45[24]), .B0(inst_cellmath__45[25]));
INVXL inst_cellmath__29_0_I2297 (.Y(N7976), .A(a_exp[1]));
INVXL inst_cellmath__29_0_I2298 (.Y(N7941), .A(a_exp[2]));
INVXL inst_cellmath__29_0_I2299 (.Y(N7950), .A(a_exp[3]));
INVXL inst_cellmath__29_0_I2300 (.Y(N7961), .A(a_exp[4]));
INVXL inst_cellmath__29_0_I2301 (.Y(N7970), .A(a_exp[5]));
INVXL inst_cellmath__29_0_I2302 (.Y(N7980), .A(a_exp[6]));
INVXL inst_cellmath__29_0_I2303 (.Y(N7945), .A(a_exp[7]));
INVXL buf1_A_I4763 (.Y(N10851), .A(N573));
INVXL buf1_A_I4764 (.Y(N7946), .A(N10851));
INVXL inst_cellmath__29_0_I2306 (.Y(N7972), .A(N7946));
AOI22XL inst_cellmath__29_0_I2308 (.Y(inst_cellmath__29[0]), .A0(N7972), .A1(N4643), .B0(N556), .B1(N7946));
AOI22XL inst_cellmath__29_0_I2309 (.Y(inst_cellmath__29[1]), .A0(N7972), .A1(N7976), .B0(N557), .B1(N7946));
AOI22XL inst_cellmath__29_0_I2310 (.Y(inst_cellmath__29[2]), .A0(N7941), .A1(N7972), .B0(N558), .B1(N7946));
AOI22XL inst_cellmath__29_0_I2311 (.Y(inst_cellmath__29[3]), .A0(N7950), .A1(N7972), .B0(N559), .B1(N7946));
AOI22XL inst_cellmath__29_0_I2312 (.Y(inst_cellmath__29[4]), .A0(N7961), .A1(N7972), .B0(N560), .B1(N7946));
AOI22XL inst_cellmath__29_0_I2313 (.Y(inst_cellmath__29[5]), .A0(N7972), .A1(N7970), .B0(N561), .B1(N7946));
AOI22XL inst_cellmath__29_0_I2314 (.Y(inst_cellmath__29[6]), .A0(N7972), .A1(N7980), .B0(N562), .B1(N7946));
AOI22XL inst_cellmath__29_0_I2315 (.Y(inst_cellmath__29[7]), .A0(N7945), .A1(N7972), .B0(N563), .B1(N7946));
NAND3XL inst_cellmath__62_0_I2317 (.Y(N8025), .A(inst_cellmath__29[6]), .B(inst_cellmath__29[7]), .C(inst_cellmath__29[5]));
NOR2XL inst_cellmath__62_0_I2318 (.Y(N8024), .A(inst_cellmath__29[0]), .B(N8025));
NAND3XL inst_cellmath__62_0_I2319 (.Y(N8021), .A(inst_cellmath__29[4]), .B(inst_cellmath__29[3]), .C(N8024));
NAND3BXL inst_cellmath__62_0_I4611 (.Y(N8015), .AN(N8021), .B(inst_cellmath__29[1]), .C(inst_cellmath__29[2]));
ADDHX1 inst_cellmath__59_0_I2332 (.CO(N8109), .S(N8088), .A(N7234), .B(inst_cellmath__29[4]));
INVXL inst_cellmath__59_0_I2333 (.Y(N8107), .A(inst_cellmath__29[7]));
ADDHX1 inst_cellmath__59_0_I11023 (.CO(N8071), .S(N17517), .A(N10734), .B(inst_cellmath__29[3]));
NOR2XL inst_cellmath__59_0_I2341 (.Y(N8053), .A(N8071), .B(N8088));
NAND2XL inst_cellmath__59_0_I2342 (.Y(N8072), .A(N8071), .B(N8088));
INVXL inst_cellmath__59_0_I2343 (.Y(N8045), .A(inst_cellmath__29[5]));
NOR2XL inst_cellmath__59_0_I2344 (.Y(N8090), .A(N8045), .B(N8109));
NAND2XL inst_cellmath__59_0_I2345 (.Y(N8110), .A(N8045), .B(N8109));
AND2XL inst_cellmath__59_0_I2346 (.Y(N8044), .A(N8045), .B(inst_cellmath__29[6]));
OR2XL inst_cellmath__59_0_I2347 (.Y(N8062), .A(N8045), .B(inst_cellmath__29[6]));
NOR2XL inst_cellmath__59_0_I2348 (.Y(N8079), .A(inst_cellmath__29[6]), .B(N8107));
NAND2XL inst_cellmath__59_0_I2349 (.Y(N8101), .A(inst_cellmath__29[6]), .B(N8107));
AOI21XL inst_cellmath__59_0_I2353 (.Y(N8066), .A0(N8110), .A1(N8053), .B0(N8090));
NAND2XL inst_cellmath__59_0_I2354 (.Y(N8083), .A(N8110), .B(N8072));
AOI21XL inst_cellmath__59_0_I2355 (.Y(N8056), .A0(N8101), .A1(N8044), .B0(N8079));
NAND2XL inst_cellmath__59_0_I2356 (.Y(N8074), .A(N8101), .B(N8062));
INVXL inst_cellmath__59_0_I2357 (.Y(N8042), .A(N8107));
OR2XL inst_cellmath__59_0_I2358 (.Y(N8058), .A(N8042), .B(N8074));
ADDHX1 inst_cellmath__59_0_I11211 (.CO(N17933), .S(N8075), .A(N7206), .B(inst_cellmath__29[0]));
XNOR2X1 inst_cellmath__59_0_I11212 (.Y(N17922), .A(N7243), .B(inst_cellmath__29[1]));
NAND2X2 inst_cellmath__59_0_I11213 (.Y(N8049), .A(N17933), .B(N17922));
NAND2X4 inst_cellmath__59_0_I11215 (.Y(N17513), .A(N8075), .B(N17525));
NOR2X2 inst_cellmath__59_0_I11216 (.Y(N8115), .A(N17933), .B(N17922));
AOI21X4 inst_cellmath__59_0_I11217 (.Y(N8087), .A0(N8049), .A1(N17513), .B0(N8115));
INVX3 inst_cellmath__59_0_I11218 (.Y(N8076), .A(N8087));
OR2XL inst_cellmath__59_0_I11021 (.Y(N17529), .A(inst_cellmath__29[1]), .B(N7243));
ADDHX1 inst_cellmath__59_0_I11022 (.CO(N17541), .S(N17535), .A(N7272), .B(inst_cellmath__29[2]));
NOR2XL inst_cellmath__59_0_I11027 (.Y(N8064), .A(N17535), .B(N17529));
NAND2XL inst_cellmath__59_0_I11028 (.Y(N8081), .A(N17535), .B(N17529));
NOR2XL inst_cellmath__59_0_I11029 (.Y(N8104), .A(N17517), .B(N17541));
NAND2XL inst_cellmath__59_0_I11030 (.Y(N8034), .A(N17541), .B(N17517));
AOI21X4 inst_cellmath__59_0_I11032 (.Y(N8078), .A0(N8064), .A1(N8034), .B0(N8104));
NAND2X1 inst_cellmath__59_0_I11033 (.Y(N8099), .A(N8034), .B(N8081));
OAI21X2 inst_cellmath__59_0_I11034 (.Y(N8068), .A0(N8099), .A1(N8087), .B0(N8078));
OAI21X2 inst_cellmath__59_0_I2361 (.Y(N8106), .A0(N8083), .A1(N8078), .B0(N8066));
NOR2XL inst_cellmath__59_0_I2362 (.Y(N8038), .A(N8083), .B(N8099));
AOI21X4 inst_cellmath__59_0_I2365 (.Y(N8048), .A0(N8038), .A1(N8076), .B0(N8106));
NAND2BXL inst_cellmath__59_0_I2366 (.Y(N8086), .AN(N8115), .B(N8049));
NAND2BXL inst_cellmath__59_0_I2367 (.Y(N8059), .AN(N8064), .B(N8081));
NAND2BXL inst_cellmath__59_0_I2368 (.Y(N8116), .AN(N8104), .B(N8034));
NAND2BXL inst_cellmath__59_0_I2369 (.Y(N8082), .AN(N8053), .B(N8072));
NAND2BXL inst_cellmath__59_0_I2370 (.Y(N8055), .AN(N8090), .B(N8110));
NAND2BXL inst_cellmath__59_0_I2371 (.Y(N8111), .AN(N8044), .B(N8062));
NAND2BXL inst_cellmath__59_0_I2372 (.Y(N8080), .AN(N8079), .B(N8101));
XNOR2X1 inst_cellmath__59_0_I2375 (.Y(inst_cellmath__59[2]), .A(N8059), .B(N8076));
XNOR2X1 inst_cellmath__59_0_I2376 (.Y(inst_cellmath__59[4]), .A(N8068), .B(N8082));
XOR2XL inst_cellmath__59_0_I2377 (.Y(inst_cellmath__59[6]), .A(N8111), .B(N8048));
XNOR2X1 inst_cellmath__59_0_I2378 (.Y(N8118), .A(N8116), .B(N8081));
XNOR2X1 inst_cellmath__59_0_I2379 (.Y(N8100), .A(N8116), .B(N8064));
MX2XL inst_cellmath__59_0_I2380 (.Y(inst_cellmath__59[3]), .A(N8100), .B(N8118), .S0(N8076));
XNOR2X1 inst_cellmath__59_0_I2381 (.Y(N8084), .A(N8055), .B(N8072));
XNOR2X1 inst_cellmath__59_0_I2382 (.Y(N8067), .A(N8055), .B(N8053));
MX2XL inst_cellmath__59_0_I2383 (.Y(inst_cellmath__59[5]), .A(N8067), .B(N8084), .S0(N8068));
XNOR2X1 inst_cellmath__59_0_I2384 (.Y(N8057), .A(N8080), .B(N8062));
XNOR2X1 inst_cellmath__59_0_I2385 (.Y(N8037), .A(N8080), .B(N8044));
MX2XL inst_cellmath__59_0_I2386 (.Y(inst_cellmath__59[7]), .A(N8057), .B(N8037), .S0(N8048));
XOR2XL inst_cellmath__59_0_I2387 (.Y(N8094), .A(N8042), .B(N8056));
NAND2XL inst_cellmath__59_0_I2388 (.Y(N8070), .A(N8074), .B(N8056));
XNOR2X1 inst_cellmath__59_0_I2389 (.Y(N8112), .A(N8042), .B(N8070));
NOR2X1 inst_cellmath__71_1_I11002 (.Y(inst_cellmath__62), .A(N8015), .B(N642));
XOR2XL inst_cellmath__71_1_I11003 (.Y(inst_cellmath__59[0]), .A(inst_cellmath__57[23]), .B(N8075));
XOR2XL inst_cellmath__71_1_I11318 (.Y(inst_cellmath__59[1]), .A(N17513), .B(N8086));
MXI2XL inst_cellmath__71_1_I11005 (.Y(N17480), .A(N8112), .B(N8094), .S0(N8048));
OAI22XL inst_cellmath__71_1_I11006 (.Y(N17489), .A0(N8058), .A1(N8048), .B0(N8042), .B1(N8056));
NAND2X2 inst_cellmath__71_1_I11007 (.Y(N17458), .A(inst_cellmath__59[2]), .B(inst_cellmath__59[5]));
NAND2X2 inst_cellmath__71_1_I11008 (.Y(N17466), .A(inst_cellmath__59[3]), .B(inst_cellmath__59[7]));
NAND2X2 inst_cellmath__71_1_I11009 (.Y(N17475), .A(inst_cellmath__59[6]), .B(inst_cellmath__59[4]));
NOR3X2 inst_cellmath__71_1_I11010 (.Y(N17485), .A(inst_cellmath__59[0]), .B(inst_cellmath__59[1]), .C(N17480));
OR4X1 inst_cellmath__71_1_I11011 (.Y(N17493), .A(N706), .B(inst_cellmath__17), .C(inst_cellmath__12), .D(inst_cellmath__63));
NOR3X4 inst_cellmath__71_1_I11012 (.Y(N17470), .A(N17458), .B(N17466), .C(N17475));
NOR2XL inst_cellmath__71_1_I11013 (.Y(N17483), .A(N17493), .B(inst_cellmath__49[5]));
NOR2XL inst_cellmath__71_1_I11014 (.Y(N17456), .A(inst_cellmath__62), .B(N17489));
NAND2X1 inst_cellmath__71_1_I11015 (.Y(N17463), .A(N17483), .B(N17456));
AOI21X4 inst_cellmath__71_1_I11016 (.Y(inst_cellmath__71), .A0(N17485), .A1(N17470), .B0(N17463));
INVX3 inst_cellmath__71_1_I4437 (.Y(N10742), .A(inst_cellmath__71));
OR3XL cynw_cm_float_add2_ieee_I4650 (.Y(N8243), .A(inst_cellmath__8), .B(inst_cellmath__4), .C(N635));
OA21X1 cynw_cm_float_add2_ieee_I4614 (.Y(N651), .A0(N634), .A1(N8243), .B0(inst_cellmath__62));
OR3XL inst_cellmath__68_0_I2409 (.Y(N8253), .A(inst_cellmath__17), .B(inst_cellmath__12), .C(inst_cellmath__63));
OR2XL inst_cellmath__68_0_I2410 (.Y(inst_cellmath__68[0]), .A(N8253), .B(N651));
NOR2XL inst_cellmath__72_0_I4615 (.Y(N8296), .A(N8253), .B(inst_cellmath__62));
INVXL inst_cellmath__72_0_I2416 (.Y(N8276), .A(inst_cellmath__59[1]));
MX2XL inst_cellmath__72_0_I11323 (.Y(x[23]), .A(inst_cellmath__59[0]), .B(inst_cellmath__68[0]), .S0(N10742));
MXI2XL inst_cellmath__72_0_I2424 (.Y(x[24]), .A(N8276), .B(N8296), .S0(N10742));
MXI2XL inst_cellmath__72_0_I2425 (.Y(x[25]), .A(inst_cellmath__59[2]), .B(N8296), .S0(N10742));
MXI2XL inst_cellmath__72_0_I2426 (.Y(x[26]), .A(inst_cellmath__59[3]), .B(N8296), .S0(N10742));
MXI2XL inst_cellmath__72_0_I11324 (.Y(x[27]), .A(inst_cellmath__59[4]), .B(N8296), .S0(N10742));
MXI2XL inst_cellmath__72_0_I2428 (.Y(x[28]), .A(inst_cellmath__59[5]), .B(N8296), .S0(N10742));
MXI2XL inst_cellmath__72_0_I2429 (.Y(x[29]), .A(inst_cellmath__59[6]), .B(N8296), .S0(N10742));
MXI2XL inst_cellmath__72_0_I2430 (.Y(x[30]), .A(inst_cellmath__59[7]), .B(N8296), .S0(N10742));
NAND3XL cynw_cm_float_add2_ieee_I2432 (.Y(N8317), .A(rm[0]), .B(rm[1]), .C(N4582));
MX2XL cynw_cm_float_add2_ieee_I2435 (.Y(N652), .A(inst_cellmath__5), .B(N7567), .S0(inst_cellmath__48));
AOI211XL inst_cellmath__70_0_I4617 (.Y(N8339), .A0(N8317), .A1(N652), .B0(inst_cellmath__8), .C0(inst_cellmath__4));
AND2XL inst_cellmath__70_0_I2438 (.Y(inst_cellmath__70), .A(N8339), .B(inst_cellmath__62));
MXI2XL inst_cellmath__73_0_I2439 (.Y(N8388), .A(inst_cellmath__70), .B(inst_cellmath__64[0]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2440 (.Y(N8417), .A(inst_cellmath__70), .B(inst_cellmath__64[1]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2441 (.Y(N8445), .A(inst_cellmath__70), .B(inst_cellmath__64[2]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2442 (.Y(N8346), .A(inst_cellmath__70), .B(inst_cellmath__64[3]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2443 (.Y(N8373), .A(inst_cellmath__70), .B(inst_cellmath__64[4]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2444 (.Y(N8400), .A(inst_cellmath__70), .B(inst_cellmath__64[5]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2445 (.Y(N8429), .A(inst_cellmath__70), .B(inst_cellmath__64[6]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2446 (.Y(N8456), .A(inst_cellmath__70), .B(inst_cellmath__64[7]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2447 (.Y(N8358), .A(inst_cellmath__70), .B(inst_cellmath__64[8]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2448 (.Y(N8384), .A(inst_cellmath__70), .B(inst_cellmath__64[9]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2449 (.Y(N8412), .A(inst_cellmath__70), .B(inst_cellmath__64[10]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2450 (.Y(N8440), .A(inst_cellmath__70), .B(inst_cellmath__64[11]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2451 (.Y(N8466), .A(inst_cellmath__70), .B(inst_cellmath__64[12]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2452 (.Y(N8368), .A(inst_cellmath__70), .B(inst_cellmath__64[13]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2453 (.Y(N8394), .A(inst_cellmath__70), .B(inst_cellmath__64[14]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2454 (.Y(N8424), .A(inst_cellmath__70), .B(inst_cellmath__64[15]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2455 (.Y(N8451), .A(inst_cellmath__70), .B(inst_cellmath__64[16]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2456 (.Y(N8353), .A(inst_cellmath__70), .B(inst_cellmath__64[17]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2457 (.Y(N8379), .A(inst_cellmath__70), .B(inst_cellmath__64[18]), .S0(inst_cellmath__63));
MX2XL inst_cellmath__73_0_I2458 (.Y(N8407), .A(inst_cellmath__70), .B(inst_cellmath__64[19]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2459 (.Y(N8435), .A(inst_cellmath__70), .B(inst_cellmath__64[20]), .S0(inst_cellmath__63));
MXI2XL inst_cellmath__73_0_I2460 (.Y(N8461), .A(inst_cellmath__70), .B(inst_cellmath__64[21]), .S0(inst_cellmath__63));
OR2XL inst_cellmath__73_0_I2461 (.Y(N8363), .A(inst_cellmath__70), .B(inst_cellmath__63));
CLKINVX6 inst_cellmath__73_0_I2486 (.Y(N8426), .A(inst_cellmath__71));
MXI2XL inst_cellmath__73_0_I2491 (.Y(x[0]), .A(inst_cellmath__57[0]), .B(N8388), .S0(N8426));
MX2XL inst_cellmath__73_0_I2492 (.Y(x[1]), .A(inst_cellmath__57[1]), .B(N8417), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2493 (.Y(x[2]), .A(inst_cellmath__57[2]), .B(N8445), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2494 (.Y(x[3]), .A(inst_cellmath__57[3]), .B(N8346), .S0(N8426));
MX2XL inst_cellmath__73_0_I2495 (.Y(x[4]), .A(inst_cellmath__57[4]), .B(N8373), .S0(N8426));
MX2XL inst_cellmath__73_0_I2496 (.Y(x[5]), .A(inst_cellmath__57[5]), .B(N8400), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2497 (.Y(x[6]), .A(inst_cellmath__57[6]), .B(N8429), .S0(N8426));
MX2XL inst_cellmath__73_0_I2498 (.Y(x[7]), .A(inst_cellmath__57[7]), .B(N8456), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2499 (.Y(x[8]), .A(inst_cellmath__57[8]), .B(N8358), .S0(N8426));
MX2XL inst_cellmath__73_0_I2500 (.Y(x[9]), .A(inst_cellmath__57[9]), .B(N8384), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2501 (.Y(x[10]), .A(inst_cellmath__57[10]), .B(N8412), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2502 (.Y(x[11]), .A(inst_cellmath__57[11]), .B(N8440), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2503 (.Y(x[12]), .A(inst_cellmath__57[12]), .B(N8466), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2504 (.Y(x[13]), .A(inst_cellmath__57[13]), .B(N8368), .S0(N8426));
MX2XL inst_cellmath__73_0_I2505 (.Y(x[14]), .A(inst_cellmath__57[14]), .B(N8394), .S0(N8426));
MX2XL inst_cellmath__73_0_I2506 (.Y(x[15]), .A(inst_cellmath__57[15]), .B(N8424), .S0(N8426));
MX2XL inst_cellmath__73_0_I2507 (.Y(x[16]), .A(inst_cellmath__57[16]), .B(N8451), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2508 (.Y(x[17]), .A(inst_cellmath__57[17]), .B(N8353), .S0(N8426));
MX2XL inst_cellmath__73_0_I2509 (.Y(x[18]), .A(inst_cellmath__57[18]), .B(N8379), .S0(N8426));
MX2XL inst_cellmath__73_0_I2510 (.Y(x[19]), .A(inst_cellmath__57[19]), .B(N8407), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2511 (.Y(x[20]), .A(inst_cellmath__57[20]), .B(N8435), .S0(N8426));
MXI2XL inst_cellmath__73_0_I2512 (.Y(x[21]), .A(inst_cellmath__57[21]), .B(N8461), .S0(N8426));
MX2XL inst_cellmath__73_0_I2513 (.Y(x[22]), .A(inst_cellmath__57[22]), .B(N8363), .S0(N8426));
assign inst_cellmath__27[3] = 1'B0;
assign inst_cellmath__27[7] = 1'B0;
assign inst_cellmath__33[0] = 1'B0;
assign inst_cellmath__33[1] = 1'B0;
assign inst_cellmath__33[2] = 1'B0;
assign inst_cellmath__33[3] = 1'B0;
assign inst_cellmath__33[4] = 1'B0;
assign inst_cellmath__33[5] = 1'B0;
assign inst_cellmath__33[6] = 1'B0;
assign inst_cellmath__33[7] = 1'B0;
assign inst_cellmath__33[8] = 1'B0;
assign inst_cellmath__33[9] = 1'B0;
assign inst_cellmath__33[10] = 1'B0;
assign inst_cellmath__33[11] = 1'B0;
assign inst_cellmath__33[12] = 1'B0;
assign inst_cellmath__33[13] = 1'B0;
assign inst_cellmath__33[14] = 1'B0;
assign inst_cellmath__33[15] = 1'B0;
assign inst_cellmath__33[16] = 1'B0;
assign inst_cellmath__33[17] = 1'B0;
assign inst_cellmath__33[18] = 1'B0;
assign inst_cellmath__33[19] = 1'B0;
assign inst_cellmath__33[20] = 1'B0;
assign inst_cellmath__33[21] = 1'B0;
assign inst_cellmath__33[22] = 1'B0;
assign inst_cellmath__33[23] = 1'B0;
assign inst_cellmath__33[25] = 1'B0;
assign inst_cellmath__33[26] = 1'B0;
assign inst_cellmath__33[30] = 1'B0;
assign inst_cellmath__33[32] = 1'B0;
assign inst_cellmath__35[0] = 1'B0;
assign inst_cellmath__36[0] = 1'B0;
assign inst_cellmath__36[1] = 1'B0;
assign inst_cellmath__36[2] = 1'B0;
assign inst_cellmath__36[3] = 1'B0;
assign inst_cellmath__36[4] = 1'B0;
assign inst_cellmath__36[5] = 1'B0;
assign inst_cellmath__36[6] = 1'B0;
assign inst_cellmath__36[7] = 1'B0;
assign inst_cellmath__36[8] = 1'B0;
assign inst_cellmath__36[9] = 1'B0;
assign inst_cellmath__36[10] = 1'B0;
assign inst_cellmath__36[11] = 1'B0;
assign inst_cellmath__36[12] = 1'B0;
assign inst_cellmath__36[13] = 1'B0;
assign inst_cellmath__36[14] = 1'B0;
assign inst_cellmath__36[15] = 1'B0;
assign inst_cellmath__36[16] = 1'B0;
assign inst_cellmath__36[17] = 1'B0;
assign inst_cellmath__36[18] = 1'B0;
assign inst_cellmath__36[19] = 1'B0;
assign inst_cellmath__36[20] = 1'B0;
assign inst_cellmath__36[21] = 1'B0;
assign inst_cellmath__36[22] = 1'B0;
assign inst_cellmath__36[23] = 1'B0;
assign inst_cellmath__36[24] = 1'B0;
assign inst_cellmath__36[25] = 1'B0;
assign inst_cellmath__36[49] = 1'B1;
assign inst_cellmath__37[25] = 1'B0;
assign inst_cellmath__37[34] = 1'B0;
assign inst_cellmath__37[35] = 1'B0;
assign inst_cellmath__37[36] = 1'B0;
assign inst_cellmath__37[37] = 1'B0;
assign inst_cellmath__37[38] = 1'B0;
assign inst_cellmath__37[39] = 1'B0;
assign inst_cellmath__37[40] = 1'B0;
assign inst_cellmath__37[41] = 1'B0;
assign inst_cellmath__37[42] = 1'B0;
assign inst_cellmath__37[43] = 1'B0;
assign inst_cellmath__37[44] = 1'B0;
assign inst_cellmath__37[45] = 1'B0;
assign inst_cellmath__37[46] = 1'B0;
assign inst_cellmath__37[47] = 1'B0;
assign inst_cellmath__37[48] = 1'B0;
assign inst_cellmath__37[49] = 1'B0;
assign inst_cellmath__39[16] = 1'B0;
assign inst_cellmath__39[24] = 1'B0;
assign inst_cellmath__45[26] = 1'B0;
assign inst_cellmath__49[2] = 1'B0;
assign inst_cellmath__49[4] = 1'B0;
assign inst_cellmath__50[0] = 1'B0;
assign inst_cellmath__59[8] = 1'B0;
assign inst_cellmath__59[9] = 1'B0;
assign inst_cellmath__64[22] = 1'B1;
assign inst_cellmath__68[1] = 1'B0;
assign inst_cellmath__68[2] = 1'B0;
assign inst_cellmath__68[3] = 1'B0;
assign inst_cellmath__68[4] = 1'B0;
assign inst_cellmath__68[5] = 1'B0;
assign inst_cellmath__68[6] = 1'B0;
assign inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  urX1QgDaqh4= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



