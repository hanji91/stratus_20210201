/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:10:45 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_0_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__5,
	inst_cellmath__7,
	inst_cellmath__10,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22;
wire [47:0] inst_cellmath__24,
	inst_cellmath__25;
wire  inst_cellmath__26,
	inst_cellmath__27,
	inst_cellmath__28;
wire [9:0] inst_cellmath__30,
	inst_cellmath__31;
wire  inst_cellmath__32,
	inst_cellmath__38,
	inst_cellmath__42,
	inst_cellmath__44;
wire [24:0] inst_cellmath__45;
wire  inst_cellmath__47;
wire [9:0] inst_cellmath__48;
wire  inst_cellmath__49;
wire N469,N1054,N1861,N2794,N2796,N2811,N2817 
	,N2827,N2830,N2832,N2836,N2838,N2842,N2848,N2852 
	,N2885,N2889,N2917,N2919,N2934,N2940,N2950,N2953 
	,N2955,N2959,N2961,N2965,N2971,N2975,N3008,N3012 
	,N3051,N3068,N3074,N3079,N3080,N3081,N3082,N3083 
	,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091 
	,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099 
	,N3100,N3101,N3103,N3105,N3106,N3107,N3108,N3109 
	,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117 
	,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125 
	,N3126,N3128,N3129,N3130,N3131,N3132,N3133,N3134 
	,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142 
	,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151 
	,N3152,N3153,N3154,N3155,N3156,N3157,N3158,N3159 
	,N3160,N3162,N3163,N3164,N3165,N3166,N3167,N3168 
	,N3169,N3171,N3172,N3174,N3175,N3176,N3177,N3178 
	,N3179,N3181,N3182,N3183,N3184,N3185,N3186,N3187 
	,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195 
	,N3196,N3197,N3198,N3200,N3201,N3202,N3203,N3205 
	,N3206,N3207,N3208,N3210,N3211,N3212,N3214,N3215 
	,N3216,N3217,N3218,N3220,N3221,N3222,N3223,N3224 
	,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232 
	,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240 
	,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248 
	,N3249,N3250,N3251,N3252,N3253,N3254,N3256,N3257 
	,N3258,N3259,N3260,N3261,N3262,N3263,N3264,N3265 
	,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3275 
	,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283 
	,N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292 
	,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300 
	,N3301,N3302,N3303,N3305,N3306,N3307,N3308,N3309 
	,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318 
	,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326 
	,N3327,N3328,N3331,N3332,N3333,N3334,N3335,N3336 
	,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344 
	,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352 
	,N3353,N3354,N3355,N3356,N3358,N3359,N3360,N3361 
	,N3362,N3364,N3365,N3366,N3367,N3368,N3369,N3370 
	,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379 
	,N3380,N3383,N3384,N3385,N3386,N3387,N3388,N3389 
	,N3390,N3391,N3392,N3393,N3394,N3396,N3397,N3398 
	,N3399,N3400,N3402,N3403,N3404,N3405,N3406,N3407 
	,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415 
	,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3424 
	,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432 
	,N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440 
	,N3441,N3442,N3443,N3444,N3446,N3447,N3448,N3449 
	,N3450,N3451,N3452,N3453,N3455,N3456,N3457,N3458 
	,N3459,N3460,N3461,N3463,N3464,N3465,N3466,N3467 
	,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475 
	,N3476,N3477,N3478,N3479,N3480,N3482,N3483,N3484 
	,N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492 
	,N3493,N3494,N3496,N3498,N3499,N3500,N3501,N3503 
	,N3504,N3505,N3506,N3507,N3508,N3510,N3512,N3513 
	,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521 
	,N3522,N3523,N3524,N3526,N3527,N3528,N3529,N3530 
	,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538 
	,N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546 
	,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554 
	,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563 
	,N3564,N3565,N3566,N3568,N3569,N3570,N3571,N3572 
	,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3581 
	,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589 
	,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597 
	,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605 
	,N3606,N3607,N3608,N3610,N3611,N3612,N3613,N3614 
	,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623 
	,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631 
	,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640 
	,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3649 
	,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657 
	,N3658,N3659,N3661,N3662,N3664,N3665,N3666,N3667 
	,N3668,N3670,N3671,N3672,N3673,N3674,N3675,N3677 
	,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685 
	,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693 
	,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701 
	,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3710 
	,N3711,N3712,N3713,N3714,N3715,N3716,N3717,N3718 
	,N3719,N3720,N3721,N3722,N3723,N3724,N3726,N3727 
	,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735 
	,N3736,N3737,N3738,N3740,N3741,N3742,N3743,N3745 
	,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753 
	,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761 
	,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3770 
	,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779 
	,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3788 
	,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796 
	,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804 
	,N3805,N3806,N3807,N3808,N3809,N3810,N3811,N3813 
	,N3814,N3815,N3816,N3817,N3818,N3819,N3821,N3822 
	,N3823,N3824,N3825,N3826,N3828,N3829,N3830,N3831 
	,N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839 
	,N3840,N3841,N3842,N3843,N3844,N3846,N3847,N3848 
	,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856 
	,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864 
	,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872 
	,N3873,N3874,N3875,N3876,N3877,N3878,N3881,N3882 
	,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890 
	,N3891,N3892,N3893,N3895,N3896,N3897,N3898,N3899 
	,N3900,N3901,N3903,N3904,N3905,N3906,N3907,N3909 
	,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917 
	,N3918,N3919,N3920,N3922,N3924,N3925,N3926,N3927 
	,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936 
	,N3937,N3938,N3940,N3941,N3942,N3943,N3944,N3945 
	,N3946,N3947,N3949,N3950,N3951,N3952,N3953,N3954 
	,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962 
	,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970 
	,N3971,N3972,N3973,N3975,N3976,N3977,N3978,N3979 
	,N3980,N3981,N3982,N3983,N3985,N3986,N3987,N3988 
	,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997 
	,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005 
	,N4006,N4007,N4008,N4010,N4011,N4012,N4013,N4014 
	,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022 
	,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031 
	,N4032,N4033,N4034,N4035,N4036,N4038,N4039,N4041 
	,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049 
	,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057 
	,N4058,N4059,N4060,N4061,N4062,N4063,N4064,N4065 
	,N4066,N4067,N4068,N4069,N4071,N4072,N4073,N4074 
	,N4075,N4077,N4078,N4079,N4080,N4081,N4082,N4084 
	,N4085,N4086,N4087,N4088,N4089,N4090,N4091,N4092 
	,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100 
	,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4109 
	,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4118 
	,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126 
	,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134 
	,N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142 
	,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150 
	,N4151,N4153,N4154,N4155,N4156,N4158,N4159,N4160 
	,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168 
	,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176 
	,N4177,N4178,N4179,N4180,N4181,N4182,N4183,N4184 
	,N4186,N4187,N4188,N4190,N4192,N4193,N4194,N4195 
	,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203 
	,N4204,N4205,N4206,N4207,N4208,N4209,N4210,N4211 
	,N4212,N4213,N4215,N4216,N4217,N4218,N4219,N4220 
	,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228 
	,N4229,N4230,N4231,N4232,N4233,N4234,N4236,N4237 
	,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245 
	,N4246,N4247,N4248,N4249,N4250,N4251,N4252,N4253 
	,N4254,N4255,N4256,N4257,N4258,N4259,N4260,N4261 
	,N4262,N4263,N4264,N4265,N4266,N4267,N4269,N4270 
	,N4271,N4272,N4273,N4274,N4275,N4278,N4279,N4280 
	,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288 
	,N4289,N4290,N4292,N4293,N4294,N4295,N4296,N4298 
	,N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306 
	,N4307,N4308,N4311,N4312,N4313,N4314,N4315,N4316 
	,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324 
	,N4325,N4326,N4327,N4328,N4329,N4330,N4331,N4332 
	,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340 
	,N4341,N4342,N4344,N4345,N4346,N4347,N4348,N4349 
	,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357 
	,N4358,N4359,N4361,N4362,N4363,N4364,N4365,N4366 
	,N4367,N4368,N4369,N4370,N4371,N4373,N4374,N4375 
	,N4376,N4377,N4378,N4379,N4380,N4382,N4383,N4384 
	,N4385,N4386,N4387,N4389,N4390,N4391,N4392,N4393 
	,N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401 
	,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409 
	,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417 
	,N4418,N4419,N4420,N4421,N4422,N4423,N4425,N4426 
	,N4427,N4428,N4430,N4431,N4432,N4433,N4435,N4436 
	,N4438,N4439,N4440,N4442,N4443,N4444,N4445,N4446 
	,N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454 
	,N4455,N4456,N4457,N4458,N4460,N4461,N4462,N4463 
	,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4473 
	,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481 
	,N4482,N4483,N4484,N4485,N4487,N4488,N4489,N4490 
	,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498 
	,N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506 
	,N4507,N4508,N4510,N4511,N4512,N4513,N4514,N4515 
	,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523 
	,N4524,N4525,N4526,N4528,N4529,N4530,N4531,N4532 
	,N4533,N4534,N4535,N4536,N4538,N4539,N4541,N4542 
	,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550 
	,N4551,N4552,N4553,N4554,N4555,N4556,N4557,N4558 
	,N4559,N4560,N4561,N4563,N4564,N4565,N4566,N4568 
	,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576 
	,N4577,N4578,N4579,N4580,N4581,N4582,N4584,N4585 
	,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4594 
	,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602 
	,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4611 
	,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619 
	,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627 
	,N4628,N4629,N4631,N4632,N4633,N4634,N4635,N4636 
	,N4637,N4638,N4639,N4640,N4641,N4643,N4644,N4645 
	,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653 
	,N4654,N4655,N4656,N4657,N4658,N4659,N4660,N4661 
	,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4670 
	,N4671,N4672,N4673,N4674,N4675,N4676,N4677,N4678 
	,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4688 
	,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696 
	,N4697,N4699,N4700,N4701,N4702,N4703,N4704,N4705 
	,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713 
	,N4714,N4715,N4716,N4717,N4718,N4720,N4721,N4722 
	,N4723,N4724,N4725,N4726,N4727,N4728,N4729,N4730 
	,N4731,N4732,N4733,N4734,N4736,N4737,N4739,N4740 
	,N4741,N4742,N4743,N4744,N4746,N4747,N4748,N4749 
	,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757 
	,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765 
	,N4766,N4767,N4768,N4769,N4770,N4771,N4772,N4773 
	,N4774,N4775,N4776,N4777,N4779,N4780,N4781,N4782 
	,N4783,N4784,N4786,N4787,N4788,N4789,N4790,N4792 
	,N4793,N4795,N4796,N4797,N4798,N4799,N4800,N4801 
	,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809 
	,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817 
	,N4818,N4819,N4821,N4822,N4823,N4824,N4825,N4826 
	,N4828,N4829,N4831,N4832,N4833,N4834,N4835,N4836 
	,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844 
	,N4845,N4846,N4847,N4848,N4849,N4850,N4851,N4852 
	,N4853,N4854,N4856,N4857,N4858,N4859,N4860,N4861 
	,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869 
	,N4870,N4871,N4872,N4873,N4874,N4876,N4877,N4878 
	,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886 
	,N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894 
	,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902 
	,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4911 
	,N4912,N4913,N4914,N4915,N4916,N4917,N4918,N4919 
	,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927 
	,N4928,N4929,N4930,N4932,N4933,N4934,N4935,N4937 
	,N4938,N4939,N4940,N4941,N4942,N4943,N4944,N4945 
	,N4946,N4947,N4948,N4949,N4950,N4952,N4953,N4954 
	,N4955,N4956,N4957,N4958,N4959,N4960,N4962,N4963 
	,N4964,N4966,N4967,N4968,N4969,N4970,N4971,N4972 
	,N4973,N4974,N4976,N4977,N4978,N4979,N4980,N4981 
	,N4982,N4983,N4984,N4985,N4986,N4988,N4989,N4990 
	,N4991,N4992,N4993,N4994,N4995,N4997,N4998,N4999 
	,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007 
	,N5009,N5010,N5011,N5012,N5014,N5016,N5017,N5018 
	,N5019,N5020,N5021,N5023,N5024,N5025,N5026,N5027 
	,N5028,N5029,N5030,N5031,N5032,N5033,N5034,N5035 
	,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043 
	,N5044,N5045,N5046,N5047,N5049,N5050,N5051,N5052 
	,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060 
	,N5061,N5062,N5064,N5065,N5066,N5067,N5068,N5069 
	,N5070,N5071,N5073,N5074,N5075,N5076,N5077,N5078 
	,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086 
	,N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094 
	,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103 
	,N5104,N5105,N5106,N5107,N5108,N5110,N5111,N5112 
	,N5113,N5114,N5115,N5116,N5117,N5119,N5120,N5121 
	,N5122,N5123,N5124,N5125,N5126,N5127,N5129,N5130 
	,N5131,N5132,N5133,N5134,N5135,N5136,N5138,N5139 
	,N5140,N5141,N5142,N5143,N5144,N5145,N7419,N7422 
	,N7424,N7425,N7428,N7429,N7430,N7432,N7433,N7435 
	,N7436,N7437,N7439,N7440,N7441,N7443,N7446,N7447 
	,N7450,N7452,N7455,N7456,N7459,N7461,N7462,N7463 
	,N7464,N7467,N7468,N7469,N7470,N7473,N7475,N7476 
	,N7478,N7479,N7481,N7482,N7484,N7485,N7486,N7490 
	,N7491,N7493,N7494,N7495,N7497,N7499,N7500,N7503 
	,N7504,N7505,N7506,N7508,N7511,N7512,N7513,N7516 
	,N7517,N7520,N7521,N7522,N7524,N7526,N7527,N7530 
	,N7532,N7534,N7537,N7538,N7540,N7543,N7545,N7546 
	,N7548,N7550,N7551,N7663,N7666,N7679,N7684,N7721 
	,N7723,N7725,N7729,N7731,N7733,N7735,N7738,N7740 
	,N7742,N7744,N7746,N7749,N7751,N7753,N7757,N7759 
	,N7761,N7763,N7848,N7849,N7852,N7854,N7857,N7859 
	,N7861,N7863,N7864,N7865,N7867,N7868,N7869,N7870 
	,N7871,N7873,N7874,N7875,N7878,N7879,N7881,N7882 
	,N7885,N7888,N7890,N7891,N7892,N7894,N7895,N7897 
	,N7898,N7899,N7900,N7902,N7903,N7904,N7907,N7908 
	,N7911,N7913,N7915,N7916,N7918,N7920,N7923,N7990 
	,N7991,N7993,N7994,N7998,N8001,N8004,N8011,N8014 
	,N8015,N8016,N8018,N8047,N8127,N8130,N8132,N8134 
	,N8136,N8138,N8140,N8157,N8173,N8176,N8178,N8181 
	,N8183,N8187,N8188,N8190,N8206,N8212,N8228,N8254 
	,N8263,N8279,N8282,N8285,N8288,N8319,N8324,N8329 
	,N8337,N8341,N8342,N8346,N8347,N8348,N8351,N8352 
	,N8354,N8360,N8361,N8363,N8368,N8371,N8373,N8374 
	,N8377,N8381,N8383,N8384,N8388,N8390,N8391,N8396 
	,N8400,N8401,N8403,N8404,N8408,N8410,N8411,N8415 
	,N8416,N8417,N8420,N8421,N8423,N8429,N8430,N8432 
	,N8434,N8439,N8440,N8442,N8446,N8447,N8450,N8452 
	,N8454,N8457,N8458,N8459,N8463,N8467,N8468,N8470 
	,N8472,N8474,N8477,N8479,N8483,N8484,N8486,N8489 
	,N8494,N8495,N8497,N8499,N8504,N8506,N8507,N8511 
	,N8512,N8515,N8519,N8522,N8524,N8525,N8526,N8529 
	,N8533,N8535,N8536,N8539,N8541,N8543,N8545,N8547 
	,N8549,N8553,N8554,N8556,N11781,N11788,N11793,N11794 
	,N11799,N11800,N11801,N11802,N11803,N11804,N11805,N11806 
	,N11807,N11813,N11821,N11829,N11836,N11840,N11847,N11854 
	,N11861,N11868,N11875,N11882,N11889,N11896,N11903,N22560 
	,N22563,N22566,N22569,N22570,N22575,N22578,N22579,N22612 
	,N22613,N22614,N22615,N22617,N22619,N22622,N22628,N22631 
	,N22634,N22637,N22638,N22641,N22643,N22646,N22677,N22678 
	,N22681,N22682,N22684,N22685,N22689,N22693,N22696,N22706 
	,N22731,N22737,N22739,N22743,N22745,N22749,N22757,N22759 
	,N22788,N22792,N22795,N22798,N22802,N22804,N22806,N22810 
	,N22815,N22816,N22818,N22819,N22846,N22848,N22852,N22854 
	,N22856,N22861,N22865,N22869,N22871,N22872,N22875,N22911 
	,N22915,N22917,N22919,N22921,N22922,N22928,N22931,N22933 
	,N22934,N22938,N22947,N22951,N22954,N22958,N22987;
NAND2XL inst_cellmath__17_0_I564 (.Y(N2796), .A(b_exp[7]), .B(b_exp[6]));
AND4XL inst_cellmath__17_0_I13953 (.Y(N2794), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL hyperpropagate_4_1_A_I5415 (.Y(N11821), .A(b_exp[0]), .B(b_exp[1]), .C(N2794));
NOR2XL hyperpropagate_4_1_A_I5416 (.Y(inst_cellmath__17), .A(N2796), .B(N11821));
NOR2XL inst_cellmath__19__2__I577 (.Y(N2817), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__19__2__I578 (.Y(N2827), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__19__2__I579 (.Y(N2838), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__19__2__I580 (.Y(N2848), .A(b_man[4]), .B(b_man[3]));
CLKINVX8 inst_cellmath__24_0_I13840 (.Y(N2811), .A(b_man[2]));
OR4X1 inst_cellmath__19__2__I13954 (.Y(N2832), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4BX1 inst_cellmath__19__2__I13957 (.Y(N2836), .AN(N2811), .B(b_man[0]), .C(N2832), .D(b_man[1]));
OR4X1 inst_cellmath__19__2__I13955 (.Y(N2842), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__19__2__I13956 (.Y(N2852), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NAND4XL inst_cellmath__19__2__I5286 (.Y(N2830), .A(N2817), .B(N2838), .C(N2827), .D(N2848));
NOR4BX1 inst_cellmath__19__2__I13958 (.Y(inst_cellmath__19), .AN(N2836), .B(N2830), .C(N2842), .D(N2852));
AND2XL cynw_cm_float_mul_ieee_I593 (.Y(inst_cellmath__21), .A(inst_cellmath__17), .B(inst_cellmath__19));
OR4X1 inst_cellmath__13__1__I13959 (.Y(N2885), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 inst_cellmath__13__1__I13960 (.Y(N2889), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL inst_cellmath__13__1__I600 (.Y(inst_cellmath__13), .A(N2885), .B(N2889));
NAND2XL inst_cellmath__10_0_I604 (.Y(N2919), .A(a_exp[7]), .B(a_exp[6]));
AND4XL inst_cellmath__10_0_I13961 (.Y(N2917), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I5417 (.Y(N11829), .A(a_exp[0]), .B(a_exp[1]), .C(N2917));
NOR2XL hyperpropagate_4_1_A_I5418 (.Y(inst_cellmath__10), .A(N2919), .B(N11829));
NOR2XL inst_cellmath__12__0__I617 (.Y(N2940), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__12__0__I618 (.Y(N2950), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__12__0__I619 (.Y(N2961), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__12__0__I620 (.Y(N2971), .A(a_man[4]), .B(a_man[3]));
CLKINVX6 inst_cellmath__12__0__I621 (.Y(N2934), .A(a_man[2]));
OR4X1 inst_cellmath__12__0__I13962 (.Y(N2955), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4BX1 inst_cellmath__12__0__I13965 (.Y(N2959), .AN(N2934), .B(a_man[0]), .C(N2955), .D(a_man[1]));
OR4X1 inst_cellmath__12__0__I13963 (.Y(N2965), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__12__0__I13964 (.Y(N2975), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NAND4XL inst_cellmath__12__0__I5288 (.Y(N2953), .A(N2940), .B(N2961), .C(N2950), .D(N2971));
NOR4BX1 inst_cellmath__12__0__I13966 (.Y(inst_cellmath__12), .AN(N2959), .B(N2953), .C(N2965), .D(N2975));
AND2XL cynw_cm_float_mul_ieee_I633 (.Y(inst_cellmath__14), .A(inst_cellmath__10), .B(inst_cellmath__12));
OR4X1 inst_cellmath__20__3__I13967 (.Y(N3008), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 inst_cellmath__20__3__I13968 (.Y(N3012), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL inst_cellmath__20__3__I640 (.Y(inst_cellmath__20), .A(N3008), .B(N3012));
NOR2BX1 cynw_cm_float_mul_ieee_I5229 (.Y(inst_cellmath__15), .AN(inst_cellmath__10), .B(inst_cellmath__12));
NOR2BX1 cynw_cm_float_mul_ieee_I5230 (.Y(inst_cellmath__22), .AN(inst_cellmath__17), .B(inst_cellmath__19));
AOI211XL cynw_cm_float_mul_ieee_I5289 (.Y(N3051), .A0(inst_cellmath__13), .A1(inst_cellmath__21), .B0(inst_cellmath__22), .C0(inst_cellmath__15));
XNOR2X1 cynw_cm_float_mul_ieee_I5234 (.Y(N11788), .A(a_sign), .B(b_sign));
NAND2BXL inst_cellmath__41_0_I654 (.Y(N3068), .AN(b_sign), .B(inst_cellmath__22));
MXI2XL inst_cellmath__41_0_I655 (.Y(N3074), .A(N3068), .B(a_sign), .S0(inst_cellmath__15));
OAI2BB1X1 inst_cellmath__31_0_I13808 (.Y(inst_cellmath__26), .A0N(inst_cellmath__20), .A1N(inst_cellmath__14), .B0(N3051));
MXI2XL inst_cellmath__41_0_I657 (.Y(x[31]), .A(N11788), .B(N3074), .S0(inst_cellmath__26));
CLKINVX6 inst_cellmath__24_0_I658 (.Y(N3346), .A(a_man[0]));
CLKINVX8 inst_cellmath__24_0_I660 (.Y(N4891), .A(a_man[1]));
CLKINVX6 inst_cellmath__24_0_I662 (.Y(N3835), .A(a_man[3]));
CLKINVX8 inst_cellmath__24_0_I664 (.Y(N3299), .A(a_man[4]));
CLKINVX8 inst_cellmath__24_0_I666 (.Y(N4845), .A(a_man[5]));
CLKINVX12 inst_cellmath__24_0_I668 (.Y(N4318), .A(a_man[6]));
CLKINVX12 inst_cellmath__24_0_I669 (.Y(N3792), .A(a_man[7]));
CLKINVX6 inst_cellmath__24_0_I670 (.Y(N3260), .A(a_man[8]));
CLKINVX8 inst_cellmath__24_0_I671 (.Y(N4801), .A(a_man[9]));
CLKINVX8 inst_cellmath__24_0_I672 (.Y(N4273), .A(a_man[10]));
CLKINVX12 inst_cellmath__24_0_I673 (.Y(N3751), .A(a_man[11]));
CLKINVX12 inst_cellmath__24_0_I674 (.Y(N3220), .A(a_man[12]));
CLKINVX8 inst_cellmath__24_0_I676 (.Y(N4758), .A(a_man[13]));
CLKINVX12 inst_cellmath__24_0_I678 (.Y(N4232), .A(a_man[14]));
CLKINVX12 inst_cellmath__24_0_I679 (.Y(N3704), .A(a_man[15]));
CLKINVX12 inst_cellmath__24_0_I680 (.Y(N3176), .A(a_man[16]));
CLKINVX16 inst_cellmath__24_0_I681 (.Y(N4715), .A(a_man[17]));
CLKINVX8 inst_cellmath__24_0_I684 (.Y(N3133), .A(a_man[20]));
CLKINVX8 inst_cellmath__24_0_I685 (.Y(N4672), .A(a_man[21]));
CLKINVX12 inst_cellmath__24_0_I686 (.Y(N4144), .A(a_man[22]));
CLKINVX12 inst_cellmath__24_0_I687 (.Y(N3620), .A(b_man[0]));
OR2X1 inst_cellmath__24_0_I689 (.Y(inst_cellmath__24[0]), .A(N3346), .B(N3620));
NOR2XL inst_cellmath__24_0_I690 (.Y(N4178), .A(N3620), .B(N4891));
NOR2XL inst_cellmath__24_0_I691 (.Y(N5084), .A(N3620), .B(N2934));
NOR2XL inst_cellmath__24_0_I692 (.Y(N3917), .A(N3620), .B(N3835));
NOR2XL inst_cellmath__24_0_I693 (.Y(N4817), .A(N3620), .B(N3299));
NOR2XL inst_cellmath__24_0_I694 (.Y(N3656), .A(N3620), .B(N4845));
NOR2XL inst_cellmath__24_0_I695 (.Y(N4558), .A(N3620), .B(N4318));
NOR2XL inst_cellmath__24_0_I696 (.Y(N3389), .A(N3620), .B(N3792));
NOR2XL inst_cellmath__24_0_I697 (.Y(N4292), .A(N3620), .B(N3260));
NOR2XL inst_cellmath__24_0_I698 (.Y(N3124), .A(N3620), .B(N4801));
NOR2XL inst_cellmath__24_0_I699 (.Y(N4031), .A(N3620), .B(N4273));
NOR2XL inst_cellmath__24_0_I700 (.Y(N4932), .A(N3620), .B(N3751));
NOR2XL inst_cellmath__24_0_I701 (.Y(N3767), .A(N3620), .B(N3220));
NOR2XL inst_cellmath__24_0_I702 (.Y(N4664), .A(N3620), .B(N4758));
NOR2XL inst_cellmath__24_0_I703 (.Y(N3505), .A(N3620), .B(N4232));
NOR2XL inst_cellmath__24_0_I704 (.Y(N4405), .A(N3620), .B(N3704));
NOR2XL inst_cellmath__24_0_I705 (.Y(N3235), .A(N3620), .B(N3176));
NOR2XL inst_cellmath__24_0_I706 (.Y(N4138), .A(N3620), .B(N4715));
CLKINVX8 inst_cellmath__24_0_I13841 (.Y(N4184), .A(a_man[18]));
NOR2XL inst_cellmath__24_0_I707 (.Y(N5042), .A(N3620), .B(N4184));
CLKINVX6 inst_cellmath__24_0_I13922 (.Y(N3666), .A(a_man[19]));
NOR2XL inst_cellmath__24_0_I708 (.Y(N3874), .A(N3620), .B(N3666));
NOR2X1 inst_cellmath__24_0_I709 (.Y(N4775), .A(N3620), .B(N3133));
NOR2XL inst_cellmath__24_0_I710 (.Y(N3612), .A(N3620), .B(N4672));
NOR2X2 inst_cellmath__24_0_I711 (.Y(N4515), .A(N3620), .B(N4144));
INVX1 inst_cellmath__24_0_I712 (.Y(N3344), .A(N3620));
CLKINVX8 inst_cellmath__24_0_I713 (.Y(N3090), .A(b_man[1]));
NOR2XL inst_cellmath__24_0_I714 (.Y(N5077), .A(N3090), .B(N3346));
NOR2XL inst_cellmath__24_0_I715 (.Y(N3907), .A(N3090), .B(N4891));
NOR2XL inst_cellmath__24_0_I716 (.Y(N4807), .A(N3090), .B(N2934));
NOR2XL inst_cellmath__24_0_I717 (.Y(N3646), .A(N3090), .B(N3835));
NOR2XL inst_cellmath__24_0_I718 (.Y(N4550), .A(N3090), .B(N3299));
NOR2XL inst_cellmath__24_0_I719 (.Y(N3378), .A(N3090), .B(N4845));
NOR2XL inst_cellmath__24_0_I720 (.Y(N4283), .A(N3090), .B(N4318));
NOR2XL inst_cellmath__24_0_I721 (.Y(N3117), .A(N3090), .B(N3792));
NOR2XL inst_cellmath__24_0_I722 (.Y(N4022), .A(N3090), .B(N3260));
NOR2XL inst_cellmath__24_0_I723 (.Y(N4923), .A(N3090), .B(N4801));
NOR2XL inst_cellmath__24_0_I724 (.Y(N3757), .A(N3090), .B(N4273));
NOR2XL inst_cellmath__24_0_I725 (.Y(N4655), .A(N3090), .B(N3751));
NOR2XL inst_cellmath__24_0_I726 (.Y(N3496), .A(N3090), .B(N3220));
NOR2XL inst_cellmath__24_0_I727 (.Y(N4396), .A(N3090), .B(N4758));
NOR2XL inst_cellmath__24_0_I728 (.Y(N3227), .A(N3090), .B(N4232));
NOR2XL inst_cellmath__24_0_I729 (.Y(N4130), .A(N3090), .B(N3704));
NOR2XL inst_cellmath__24_0_I730 (.Y(N5035), .A(N3090), .B(N3176));
NOR2XL inst_cellmath__24_0_I731 (.Y(N3865), .A(N3090), .B(N4715));
NOR2XL inst_cellmath__24_0_I732 (.Y(N4766), .A(N3090), .B(N4184));
NOR2X2 inst_cellmath__24_0_I733 (.Y(N3601), .A(N3090), .B(N3666));
NOR2XL inst_cellmath__24_0_I734 (.Y(N4506), .A(N3090), .B(N3133));
NOR2X1 inst_cellmath__24_0_I735 (.Y(N3335), .A(N4672), .B(N3090));
NOR2X1 inst_cellmath__24_0_I736 (.Y(N4238), .A(N3090), .B(N4144));
INVX1 inst_cellmath__24_0_I737 (.Y(N5142), .A(N3090));
NOR2XL inst_cellmath__24_0_I740 (.Y(N4798), .A(N2811), .B(N3346));
NOR2XL inst_cellmath__24_0_I741 (.Y(N3637), .A(N2811), .B(N4891));
NOR2XL inst_cellmath__24_0_I742 (.Y(N4541), .A(N2811), .B(N2934));
NOR2XL inst_cellmath__24_0_I743 (.Y(N3367), .A(N2811), .B(N3835));
NOR2XL inst_cellmath__24_0_I744 (.Y(N4272), .A(N2811), .B(N3299));
NOR2XL inst_cellmath__24_0_I745 (.Y(N3108), .A(N2811), .B(N4845));
NOR2XL inst_cellmath__24_0_I746 (.Y(N4013), .A(N2811), .B(N4318));
NOR2XL inst_cellmath__24_0_I747 (.Y(N4914), .A(N2811), .B(N3792));
NOR2XL inst_cellmath__24_0_I748 (.Y(N3748), .A(N2811), .B(N3260));
NOR2XL inst_cellmath__24_0_I749 (.Y(N4645), .A(N2811), .B(N4801));
NOR2XL inst_cellmath__24_0_I750 (.Y(N3486), .A(N2811), .B(N4273));
NOR2XL inst_cellmath__24_0_I751 (.Y(N4385), .A(N2811), .B(N3751));
NOR2XL inst_cellmath__24_0_I752 (.Y(N3216), .A(N2811), .B(N3220));
NOR2XL inst_cellmath__24_0_I753 (.Y(N4122), .A(N2811), .B(N4758));
NOR2XL inst_cellmath__24_0_I754 (.Y(N5026), .A(N2811), .B(N4232));
NOR2XL inst_cellmath__24_0_I755 (.Y(N3857), .A(N3704), .B(N2811));
NOR2XL inst_cellmath__24_0_I756 (.Y(N4757), .A(N2811), .B(N3176));
NOR2XL inst_cellmath__24_0_I757 (.Y(N3592), .A(N4715), .B(N2811));
NOR2X2 inst_cellmath__24_0_I13842 (.Y(N4498), .A(N4184), .B(N2811));
NOR2X1 inst_cellmath__24_0_I759 (.Y(N3323), .A(N2811), .B(N3666));
NOR2X2 inst_cellmath__24_0_I760 (.Y(N4228), .A(N2811), .B(N3133));
NOR2X2 inst_cellmath__24_0_I761 (.Y(N5132), .A(N4672), .B(N2811));
NOR2X2 inst_cellmath__24_0_I762 (.Y(N3968), .A(N4144), .B(N2811));
INVX1 inst_cellmath__24_0_I763 (.Y(N4868), .A(N2811));
CLKINVX16 inst_cellmath__24_0_I764 (.Y(N3655), .A(b_man[3]));
NOR2XL inst_cellmath__24_0_I766 (.Y(N4531), .A(N3655), .B(N3346));
NOR2XL inst_cellmath__24_0_I767 (.Y(N3358), .A(N3655), .B(N4891));
NOR2XL inst_cellmath__24_0_I768 (.Y(N4260), .A(N3655), .B(N2934));
NOR2XL inst_cellmath__24_0_I769 (.Y(N3097), .A(N3655), .B(N3835));
NOR2XL inst_cellmath__24_0_I770 (.Y(N4003), .A(N3655), .B(N3299));
NOR2XL inst_cellmath__24_0_I771 (.Y(N4903), .A(N4845), .B(N3655));
NOR2XL inst_cellmath__24_0_I772 (.Y(N3738), .A(N3655), .B(N4318));
NOR2XL inst_cellmath__24_0_I773 (.Y(N4636), .A(N3655), .B(N3792));
NOR2XL inst_cellmath__24_0_I774 (.Y(N3475), .A(N3655), .B(N3260));
NOR2XL inst_cellmath__24_0_I775 (.Y(N4374), .A(N3655), .B(N4801));
NOR2XL inst_cellmath__24_0_I776 (.Y(N3206), .A(N3655), .B(N4273));
NOR2XL inst_cellmath__24_0_I777 (.Y(N4111), .A(N3655), .B(N3751));
NOR2XL inst_cellmath__24_0_I778 (.Y(N5016), .A(N3655), .B(N3220));
NOR2XL inst_cellmath__24_0_I779 (.Y(N3847), .A(N3655), .B(N4758));
NOR2X1 inst_cellmath__24_0_I780 (.Y(N4748), .A(N3655), .B(N4232));
NOR2XL inst_cellmath__24_0_I781 (.Y(N3582), .A(N3655), .B(N3704));
NOR2X1 inst_cellmath__24_0_I782 (.Y(N4488), .A(N3655), .B(N3176));
NOR2X2 inst_cellmath__24_0_I783 (.Y(N3314), .A(N3655), .B(N4715));
NOR2X1 inst_cellmath__24_0_I784 (.Y(N4217), .A(N3655), .B(N4184));
NOR2X1 inst_cellmath__24_0_I785 (.Y(N5120), .A(N3655), .B(N3666));
NOR2X1 inst_cellmath__24_0_I786 (.Y(N3958), .A(N3655), .B(N3133));
NOR2XL inst_cellmath__24_0_I787 (.Y(N4859), .A(N3655), .B(N4672));
NOR2X1 inst_cellmath__24_0_I788 (.Y(N3695), .A(N4144), .B(N3655));
INVXL inst_cellmath__24_0_I789 (.Y(N4596), .A(N3655));
CLKINVX8 inst_cellmath__24_0_I790 (.Y(N4737), .A(b_man[4]));
INVX8 inst_cellmath__24_0_I5122 (.Y(N11793), .A(N4737));
INVX12 inst_cellmath__24_0_I5123 (.Y(N11794), .A(N11793));
NOR2XL inst_cellmath__24_0_I793 (.Y(N4252), .A(N11794), .B(N3346));
NOR2XL inst_cellmath__24_0_I794 (.Y(N3087), .A(N11794), .B(N4891));
NOR2XL inst_cellmath__24_0_I795 (.Y(N3993), .A(N11794), .B(N2934));
NOR2XL inst_cellmath__24_0_I796 (.Y(N4895), .A(N11794), .B(N3835));
NOR2XL inst_cellmath__24_0_I797 (.Y(N3729), .A(N3299), .B(N11794));
NOR2XL inst_cellmath__24_0_I798 (.Y(N4627), .A(N11794), .B(N4845));
NOR2XL inst_cellmath__24_0_I799 (.Y(N3466), .A(N11794), .B(N4318));
NOR2XL inst_cellmath__24_0_I800 (.Y(N4365), .A(N11794), .B(N3792));
NOR2XL inst_cellmath__24_0_I801 (.Y(N3196), .A(N11794), .B(N3260));
NOR2XL inst_cellmath__24_0_I802 (.Y(N4102), .A(N11794), .B(N4801));
NOR2XL inst_cellmath__24_0_I803 (.Y(N5005), .A(N11794), .B(N4273));
NOR2XL inst_cellmath__24_0_I804 (.Y(N3838), .A(N11794), .B(N3751));
NOR2XL inst_cellmath__24_0_I805 (.Y(N4736), .A(N3220), .B(N11794));
NOR2X1 inst_cellmath__24_0_I806 (.Y(N3573), .A(N4758), .B(N11794));
NOR2XL inst_cellmath__24_0_I807 (.Y(N4479), .A(N11794), .B(N4232));
NOR2XL inst_cellmath__24_0_I808 (.Y(N3303), .A(N4737), .B(N3704));
NOR2X1 inst_cellmath__24_0_I809 (.Y(N4208), .A(N3176), .B(N4737));
NOR2X4 inst_cellmath__24_0_I810 (.Y(N5111), .A(N4715), .B(N11794));
NOR2X2 inst_cellmath__24_0_I811 (.Y(N3947), .A(N4184), .B(N4737));
NOR2X1 inst_cellmath__24_0_I812 (.Y(N4848), .A(N4737), .B(N3666));
NOR2X1 inst_cellmath__24_0_I813 (.Y(N3684), .A(N4737), .B(N3133));
NOR2X4 inst_cellmath__24_0_I814 (.Y(N4587), .A(N4672), .B(N11794));
NOR2X4 inst_cellmath__24_0_I815 (.Y(N3420), .A(N4144), .B(N11794));
INVXL inst_cellmath__24_0_I816 (.Y(N4320), .A(N11794));
CLKINVX8 inst_cellmath__24_0_I13923 (.Y(N3766), .A(b_man[5]));
NOR2XL inst_cellmath__24_0_I820 (.Y(N3985), .A(N3766), .B(N3346));
NOR2XL inst_cellmath__24_0_I821 (.Y(N4886), .A(N3766), .B(N4891));
NOR2XL inst_cellmath__24_0_I822 (.Y(N3720), .A(N3766), .B(N2934));
NOR2XL inst_cellmath__24_0_I823 (.Y(N4619), .A(N3766), .B(N3835));
NOR2XL inst_cellmath__24_0_I824 (.Y(N3458), .A(N3766), .B(N3299));
NOR2XL inst_cellmath__24_0_I825 (.Y(N4354), .A(N3766), .B(N4845));
NOR2XL inst_cellmath__24_0_I826 (.Y(N3188), .A(N3766), .B(N4318));
NOR2XL inst_cellmath__24_0_I827 (.Y(N4094), .A(N3766), .B(N3792));
NOR2XL inst_cellmath__24_0_I4992 (.Y(N11781), .A(N3766), .B(N3260));
NOR2XL inst_cellmath__24_0_I829 (.Y(N3829), .A(N3766), .B(N4801));
NOR2XL inst_cellmath__24_0_I830 (.Y(N4727), .A(N3766), .B(N4273));
NOR2XL inst_cellmath__24_0_I831 (.Y(N3563), .A(N3766), .B(N3751));
NOR2XL inst_cellmath__24_0_I832 (.Y(N4468), .A(N3766), .B(N3220));
NOR2XL inst_cellmath__24_0_I833 (.Y(N3294), .A(N4758), .B(N3766));
NOR2X1 inst_cellmath__24_0_I834 (.Y(N4199), .A(N3766), .B(N4232));
NOR2X2 inst_cellmath__24_0_I835 (.Y(N5104), .A(N3704), .B(N3766));
NOR2X1 inst_cellmath__24_0_I836 (.Y(N3938), .A(N3766), .B(N3176));
NOR2X4 inst_cellmath__24_0_I837 (.Y(N4839), .A(N3766), .B(N4715));
NOR2X2 inst_cellmath__24_0_I838 (.Y(N3677), .A(N3766), .B(N4184));
NOR2X1 inst_cellmath__24_0_I13924 (.Y(N4577), .A(N3666), .B(N3766));
NOR2X1 inst_cellmath__24_0_I840 (.Y(N3410), .A(N3766), .B(N3133));
NOR2X1 inst_cellmath__24_0_I841 (.Y(N4312), .A(N3766), .B(N4672));
NOR2XL inst_cellmath__24_0_I842 (.Y(N3146), .A(N3766), .B(N4144));
INVXL inst_cellmath__24_0_I843 (.Y(N4052), .A(N3766));
CLKINVX8 inst_cellmath__24_0_I844 (.Y(N4851), .A(b_man[6]));
NOR2XL inst_cellmath__24_0_I846 (.Y(N3711), .A(N4851), .B(N3346));
NOR2XL inst_cellmath__24_0_I847 (.Y(N4609), .A(N4851), .B(N4891));
NOR2XL inst_cellmath__24_0_I848 (.Y(N3444), .A(N4851), .B(N2934));
NOR2XL inst_cellmath__24_0_I849 (.Y(N4345), .A(N4851), .B(N3835));
NOR2XL inst_cellmath__24_0_I850 (.Y(N3179), .A(N4851), .B(N3299));
NOR2XL inst_cellmath__24_0_I851 (.Y(N4082), .A(N4851), .B(N4845));
NOR2XL inst_cellmath__24_0_I852 (.Y(N4989), .A(N4851), .B(N4318));
NOR2XL inst_cellmath__24_0_I853 (.Y(N3819), .A(N4851), .B(N3792));
NOR2XL inst_cellmath__24_0_I854 (.Y(N4718), .A(N4851), .B(N3260));
NOR2XL inst_cellmath__24_0_I855 (.Y(N3554), .A(N4851), .B(N4801));
NOR2XL inst_cellmath__24_0_I856 (.Y(N4458), .A(N4851), .B(N4273));
NOR2XL inst_cellmath__24_0_I857 (.Y(N3287), .A(N3751), .B(N4851));
NOR2X1 inst_cellmath__24_0_I858 (.Y(N4190), .A(N3220), .B(N4851));
NOR2X1 inst_cellmath__24_0_I859 (.Y(N5094), .A(N4851), .B(N4758));
NOR2X4 inst_cellmath__24_0_I860 (.Y(N3930), .A(N4232), .B(N4851));
NOR2X1 inst_cellmath__24_0_I861 (.Y(N4829), .A(N3704), .B(N4851));
NOR2X2 inst_cellmath__24_0_I862 (.Y(N3668), .A(N3176), .B(N4851));
NOR2X2 inst_cellmath__24_0_I863 (.Y(N4570), .A(N4715), .B(N4851));
NOR2X1 inst_cellmath__24_0_I864 (.Y(N3400), .A(N4184), .B(N4851));
NOR2XL inst_cellmath__24_0_I865 (.Y(N4302), .A(N4851), .B(N3666));
NOR2X1 inst_cellmath__24_0_I866 (.Y(N3138), .A(N3133), .B(N4851));
NOR2X1 inst_cellmath__24_0_I867 (.Y(N4043), .A(N4851), .B(N4672));
NOR2XL inst_cellmath__24_0_I868 (.Y(N4942), .A(N4851), .B(N4144));
INVXL inst_cellmath__24_0_I869 (.Y(N3781), .A(N4851));
CLKINVX12 inst_cellmath__24_0_I870 (.Y(N4324), .A(b_man[7]));
NOR2XL inst_cellmath__24_0_I872 (.Y(N3435), .A(N4324), .B(N3346));
NOR2XL inst_cellmath__24_0_I873 (.Y(N4335), .A(N4324), .B(N4891));
NOR2XL inst_cellmath__24_0_I874 (.Y(N3168), .A(N4324), .B(N2934));
NOR2XL inst_cellmath__24_0_I875 (.Y(N4073), .A(N4324), .B(N3835));
NOR2XL inst_cellmath__24_0_I876 (.Y(N4980), .A(N4324), .B(N3299));
NOR2XL inst_cellmath__24_0_I877 (.Y(N3811), .A(N4324), .B(N4845));
NOR2XL inst_cellmath__24_0_I878 (.Y(N4709), .A(N4324), .B(N4318));
NOR2XL inst_cellmath__24_0_I879 (.Y(N3547), .A(N4324), .B(N3792));
NOR2XL inst_cellmath__24_0_I880 (.Y(N4451), .A(N4324), .B(N3260));
NOR2XL inst_cellmath__24_0_I881 (.Y(N3277), .A(N4324), .B(N4801));
NOR2XL inst_cellmath__24_0_I882 (.Y(N4181), .A(N4324), .B(N4273));
NOR2X1 inst_cellmath__24_0_I883 (.Y(N5087), .A(N3751), .B(N4324));
NOR2XL inst_cellmath__24_0_I884 (.Y(N3920), .A(N4324), .B(N3220));
NOR2XL inst_cellmath__24_0_I885 (.Y(N4822), .A(N4324), .B(N4758));
NOR2X1 inst_cellmath__24_0_I886 (.Y(N3659), .A(N4324), .B(N4232));
NOR2X1 inst_cellmath__24_0_I887 (.Y(N4561), .A(N4324), .B(N3704));
NOR2X2 inst_cellmath__24_0_I888 (.Y(N3394), .A(N4324), .B(N3176));
NOR2XL inst_cellmath__24_0_I889 (.Y(N4296), .A(N4324), .B(N4715));
NOR2XL inst_cellmath__24_0_I890 (.Y(N3130), .A(N4324), .B(N4184));
NOR2XL inst_cellmath__24_0_I891 (.Y(N4036), .A(N4324), .B(N3666));
NOR2XL inst_cellmath__24_0_I892 (.Y(N4935), .A(N4324), .B(N3133));
NOR2XL inst_cellmath__24_0_I893 (.Y(N3774), .A(N4324), .B(N4672));
NOR2XL inst_cellmath__24_0_I894 (.Y(N4668), .A(N4324), .B(N4144));
INVXL inst_cellmath__24_0_I895 (.Y(N3508), .A(N4324));
CLKINVX12 inst_cellmath__24_0_I896 (.Y(N3798), .A(b_man[8]));
NOR2XL inst_cellmath__24_0_I898 (.Y(N3160), .A(N3798), .B(N3346));
NOR2XL inst_cellmath__24_0_I899 (.Y(N4064), .A(N3798), .B(N4891));
NOR2XL inst_cellmath__24_0_I900 (.Y(N4970), .A(N3798), .B(N2934));
NOR2XL inst_cellmath__24_0_I901 (.Y(N3803), .A(N3798), .B(N3835));
NOR2XL inst_cellmath__24_0_I902 (.Y(N4701), .A(N3798), .B(N3299));
NOR2XL inst_cellmath__24_0_I903 (.Y(N3539), .A(N3798), .B(N4845));
NOR2XL inst_cellmath__24_0_I904 (.Y(N4443), .A(N3798), .B(N4318));
NOR2XL inst_cellmath__24_0_I905 (.Y(N3269), .A(N3798), .B(N3792));
NOR2XL inst_cellmath__24_0_I906 (.Y(N4173), .A(N3798), .B(N3260));
NOR2XL inst_cellmath__24_0_I907 (.Y(N5079), .A(N3798), .B(N4801));
NOR2X1 inst_cellmath__24_0_I908 (.Y(N3911), .A(N4273), .B(N3798));
NOR2XL inst_cellmath__24_0_I909 (.Y(N4811), .A(N3798), .B(N3751));
NOR2X2 inst_cellmath__24_0_I910 (.Y(N3649), .A(N3220), .B(N3798));
NOR2X2 inst_cellmath__24_0_I911 (.Y(N4553), .A(N3798), .B(N4758));
NOR2X1 inst_cellmath__24_0_I912 (.Y(N3384), .A(N4232), .B(N3798));
NOR2X1 inst_cellmath__24_0_I913 (.Y(N4285), .A(N3704), .B(N3798));
NOR2X2 inst_cellmath__24_0_I914 (.Y(N3120), .A(N3176), .B(N3798));
NOR2X2 inst_cellmath__24_0_I915 (.Y(N4026), .A(N3798), .B(N4715));
NOR2X1 inst_cellmath__24_0_I916 (.Y(N4927), .A(N3798), .B(N4184));
NOR2XL inst_cellmath__24_0_I917 (.Y(N3760), .A(N3798), .B(N3666));
NOR2XL inst_cellmath__24_0_I918 (.Y(N4660), .A(N3133), .B(N3798));
NOR2XL inst_cellmath__24_0_I919 (.Y(N3501), .A(N3798), .B(N4672));
NOR2XL inst_cellmath__24_0_I920 (.Y(N4400), .A(N3798), .B(N4144));
INVXL inst_cellmath__24_0_I921 (.Y(N3231), .A(N3798));
CLKINVX8 inst_cellmath__24_0_I922 (.Y(N4887), .A(b_man[9]));
NOR2XL inst_cellmath__24_0_I924 (.Y(N4960), .A(N4887), .B(N3346));
NOR2XL inst_cellmath__24_0_I925 (.Y(N3794), .A(N4887), .B(N4891));
NOR2XL inst_cellmath__24_0_I926 (.Y(N4692), .A(N4887), .B(N2934));
NOR2XL inst_cellmath__24_0_I927 (.Y(N3533), .A(N4887), .B(N3835));
NOR2XL inst_cellmath__24_0_I928 (.Y(N4432), .A(N4887), .B(N3299));
NOR2XL inst_cellmath__24_0_I929 (.Y(N3261), .A(N4887), .B(N4845));
NOR2XL inst_cellmath__24_0_I930 (.Y(N4165), .A(N4318), .B(N4887));
NOR2XL inst_cellmath__24_0_I931 (.Y(N5069), .A(N4887), .B(N3792));
NOR2XL inst_cellmath__24_0_I932 (.Y(N3900), .A(N4887), .B(N3260));
NOR2XL inst_cellmath__24_0_I933 (.Y(N4803), .A(N4887), .B(N4801));
NOR2XL inst_cellmath__24_0_I934 (.Y(N3639), .A(N4887), .B(N4273));
NOR2X2 inst_cellmath__24_0_I935 (.Y(N4545), .A(N3751), .B(N4887));
NOR2X2 inst_cellmath__24_0_I936 (.Y(N3372), .A(N3220), .B(N4887));
NOR2X2 inst_cellmath__24_0_I937 (.Y(N4275), .A(N4758), .B(N4887));
NOR2X2 inst_cellmath__24_0_I938 (.Y(N3112), .A(N4232), .B(N4887));
NOR2X2 inst_cellmath__24_0_I939 (.Y(N4017), .A(N3704), .B(N4887));
NOR2X2 inst_cellmath__24_0_I940 (.Y(N4916), .A(N3176), .B(N4887));
NOR2X1 inst_cellmath__24_0_I941 (.Y(N3752), .A(N4715), .B(N4887));
NOR2XL inst_cellmath__24_0_I942 (.Y(N4650), .A(N4887), .B(N4184));
NOR2XL inst_cellmath__24_0_I943 (.Y(N3490), .A(N4887), .B(N3666));
NOR2XL inst_cellmath__24_0_I944 (.Y(N4389), .A(N4887), .B(N3133));
NOR2XL inst_cellmath__24_0_I945 (.Y(N3223), .A(N4887), .B(N4672));
NOR2XL inst_cellmath__24_0_I946 (.Y(N4125), .A(N4887), .B(N4144));
INVXL inst_cellmath__24_0_I947 (.Y(N5029), .A(N4887));
CLKINVX8 inst_cellmath__24_0_I948 (.Y(N3906), .A(b_man[10]));
NOR2XL inst_cellmath__24_0_I950 (.Y(N4683), .A(N3906), .B(N3346));
NOR2XL inst_cellmath__24_0_I951 (.Y(N3523), .A(N3906), .B(N4891));
NOR2XL inst_cellmath__24_0_I952 (.Y(N4422), .A(N3906), .B(N2934));
NOR2XL inst_cellmath__24_0_I953 (.Y(N3252), .A(N3906), .B(N3835));
NOR2XL inst_cellmath__24_0_I954 (.Y(N4156), .A(N3906), .B(N3299));
NOR2XL inst_cellmath__24_0_I955 (.Y(N5061), .A(N3906), .B(N4845));
NOR2XL inst_cellmath__24_0_I956 (.Y(N3891), .A(N3906), .B(N4318));
NOR2XL inst_cellmath__24_0_I957 (.Y(N4793), .A(N3906), .B(N3792));
NOR2X1 inst_cellmath__24_0_I958 (.Y(N3629), .A(N3906), .B(N3260));
NOR2XL inst_cellmath__24_0_I959 (.Y(N4534), .A(N3906), .B(N4801));
NOR2XL inst_cellmath__24_0_I960 (.Y(N3362), .A(N3906), .B(N4273));
NOR2X1 inst_cellmath__24_0_I961 (.Y(N4263), .A(N3751), .B(N3906));
NOR2X2 inst_cellmath__24_0_I962 (.Y(N3100), .A(N3906), .B(N3220));
NOR2X1 inst_cellmath__24_0_I963 (.Y(N4008), .A(N3906), .B(N4758));
NOR2X1 inst_cellmath__24_0_I964 (.Y(N4905), .A(N3906), .B(N4232));
NOR2X1 inst_cellmath__24_0_I965 (.Y(N3742), .A(N3906), .B(N3704));
NOR2XL inst_cellmath__24_0_I966 (.Y(N4640), .A(N3906), .B(N3176));
NOR2XL inst_cellmath__24_0_I967 (.Y(N3478), .A(N3906), .B(N4715));
NOR2XL inst_cellmath__24_0_I968 (.Y(N4378), .A(N3906), .B(N4184));
NOR2XL inst_cellmath__24_0_I969 (.Y(N3212), .A(N3906), .B(N3666));
NOR2XL inst_cellmath__24_0_I970 (.Y(N4114), .A(N3906), .B(N3133));
NOR2XL inst_cellmath__24_0_I971 (.Y(N5019), .A(N3906), .B(N4672));
NOR2XL inst_cellmath__24_0_I972 (.Y(N3852), .A(N3906), .B(N4144));
INVXL inst_cellmath__24_0_I973 (.Y(N4751), .A(N3906));
CLKINVX8 inst_cellmath__24_0_I974 (.Y(N3376), .A(b_man[11]));
NOR2XL inst_cellmath__24_0_I975 (.Y(N4414), .A(N3376), .B(N3346));
NOR2XL inst_cellmath__24_0_I976 (.Y(N3242), .A(N3376), .B(N4891));
NOR2XL inst_cellmath__24_0_I977 (.Y(N4145), .A(N3376), .B(N2934));
NOR2XL inst_cellmath__24_0_I978 (.Y(N5052), .A(N3376), .B(N3835));
NOR2XL inst_cellmath__24_0_I979 (.Y(N3882), .A(N3376), .B(N3299));
NOR2XL inst_cellmath__24_0_I980 (.Y(N4782), .A(N3376), .B(N4845));
NOR2XL inst_cellmath__24_0_I981 (.Y(N3623), .A(N3376), .B(N4318));
NOR2XL inst_cellmath__24_0_I982 (.Y(N4522), .A(N3376), .B(N3792));
NOR2XL inst_cellmath__24_0_I983 (.Y(N3352), .A(N3376), .B(N3260));
NOR2XL inst_cellmath__24_0_I984 (.Y(N4255), .A(N3376), .B(N4801));
NOR2X2 inst_cellmath__24_0_I985 (.Y(N3091), .A(N4273), .B(N3376));
NOR2XL inst_cellmath__24_0_I986 (.Y(N3996), .A(N3751), .B(N3376));
NOR2X2 inst_cellmath__24_0_I987 (.Y(N4898), .A(N3220), .B(N3376));
NOR2X2 inst_cellmath__24_0_I988 (.Y(N3732), .A(N4758), .B(N3376));
NOR2X1 inst_cellmath__24_0_I989 (.Y(N4633), .A(N3376), .B(N4232));
NOR2XL inst_cellmath__24_0_I990 (.Y(N3469), .A(N3704), .B(N3376));
NOR2XL inst_cellmath__24_0_I991 (.Y(N4368), .A(N3376), .B(N3176));
NOR2XL inst_cellmath__24_0_I992 (.Y(N3202), .A(N3376), .B(N4715));
NOR2XL inst_cellmath__24_0_I993 (.Y(N4105), .A(N3376), .B(N4184));
NOR2XL inst_cellmath__24_0_I994 (.Y(N5009), .A(N3376), .B(N3666));
NOR2XL inst_cellmath__24_0_I995 (.Y(N3843), .A(N3376), .B(N3133));
NOR2XL inst_cellmath__24_0_I996 (.Y(N4741), .A(N3376), .B(N4672));
NOR2XL inst_cellmath__24_0_I997 (.Y(N3576), .A(N3376), .B(N4144));
INVXL inst_cellmath__24_0_I998 (.Y(N4484), .A(N3376));
CLKINVX8 inst_cellmath__24_0_I999 (.Y(N4922), .A(b_man[12]));
NOR2XL inst_cellmath__24_0_I1002 (.Y(N4137), .A(N4922), .B(N3346));
NOR2XL inst_cellmath__24_0_I1003 (.Y(N5044), .A(N4922), .B(N4891));
NOR2XL inst_cellmath__24_0_I1004 (.Y(N3873), .A(N4922), .B(N2934));
NOR2XL inst_cellmath__24_0_I1005 (.Y(N4774), .A(N4922), .B(N3835));
NOR2XL inst_cellmath__24_0_I1006 (.Y(N3614), .A(N4922), .B(N3299));
NOR2XL inst_cellmath__24_0_I1007 (.Y(N4514), .A(N4922), .B(N4845));
NOR2XL inst_cellmath__24_0_I1008 (.Y(N3343), .A(N4922), .B(N4318));
NOR2X1 inst_cellmath__24_0_I1009 (.Y(N4248), .A(N3792), .B(N4922));
NOR2X1 inst_cellmath__24_0_I1010 (.Y(N3082), .A(N3260), .B(N4922));
NOR2X2 inst_cellmath__24_0_I1011 (.Y(N3988), .A(N4801), .B(N4922));
NOR2X1 inst_cellmath__24_0_I1012 (.Y(N4890), .A(N4922), .B(N4273));
NOR2X1 inst_cellmath__24_0_I1013 (.Y(N3724), .A(N3751), .B(N4922));
NOR2X2 inst_cellmath__24_0_I1014 (.Y(N4622), .A(N4922), .B(N3220));
NOR2XL inst_cellmath__24_0_I1015 (.Y(N3461), .A(N4922), .B(N4758));
NOR2X1 inst_cellmath__24_0_I1016 (.Y(N4359), .A(N4922), .B(N4232));
NOR2XL inst_cellmath__24_0_I1017 (.Y(N3191), .A(N3704), .B(N4922));
NOR2X1 inst_cellmath__24_0_I1018 (.Y(N4098), .A(N3176), .B(N4922));
NOR2XL inst_cellmath__24_0_I1019 (.Y(N5001), .A(N4922), .B(N4715));
NOR2XL inst_cellmath__24_0_I1020 (.Y(N3832), .A(N4922), .B(N4184));
NOR2XL inst_cellmath__24_0_I1021 (.Y(N4731), .A(N4922), .B(N3666));
NOR2XL inst_cellmath__24_0_I1022 (.Y(N3569), .A(N4922), .B(N3133));
NOR2XL inst_cellmath__24_0_I1023 (.Y(N4476), .A(N4922), .B(N4672));
NOR2XL inst_cellmath__24_0_I1024 (.Y(N3298), .A(N4922), .B(N4144));
INVXL inst_cellmath__24_0_I1025 (.Y(N4203), .A(N4922));
CLKINVX6 inst_cellmath__24_0_I1026 (.Y(N4395), .A(b_man[13]));
NOR2XL inst_cellmath__24_0_I1028 (.Y(N3864), .A(N4395), .B(N3346));
NOR2XL inst_cellmath__24_0_I1029 (.Y(N4765), .A(N4395), .B(N4891));
NOR2XL inst_cellmath__24_0_I1030 (.Y(N3604), .A(N4395), .B(N2934));
NOR2XL inst_cellmath__24_0_I1031 (.Y(N4505), .A(N4395), .B(N3835));
NOR2XL inst_cellmath__24_0_I1032 (.Y(N3334), .A(N4395), .B(N3299));
NOR2XL inst_cellmath__24_0_I1033 (.Y(N4241), .A(N4395), .B(N4845));
NOR2X1 inst_cellmath__24_0_I1034 (.Y(N5141), .A(N4318), .B(N4395));
NOR2X1 inst_cellmath__24_0_I1035 (.Y(N3979), .A(N3792), .B(N4395));
NOR2X1 inst_cellmath__24_0_I1036 (.Y(N4880), .A(N3260), .B(N4395));
NOR2XL inst_cellmath__24_0_I1037 (.Y(N3714), .A(N4395), .B(N4801));
NOR2X1 inst_cellmath__24_0_I1038 (.Y(N4613), .A(N4395), .B(N4273));
NOR2X1 inst_cellmath__24_0_I1039 (.Y(N3451), .A(N4395), .B(N3751));
NOR2X2 inst_cellmath__24_0_I1040 (.Y(N4348), .A(N4395), .B(N3220));
NOR2X1 inst_cellmath__24_0_I1041 (.Y(N3183), .A(N4395), .B(N4758));
NOR2XL inst_cellmath__24_0_I1042 (.Y(N4088), .A(N4395), .B(N4232));
NOR2XL inst_cellmath__24_0_I1043 (.Y(N4993), .A(N4395), .B(N3704));
NOR2XL inst_cellmath__24_0_I1044 (.Y(N3824), .A(N4395), .B(N3176));
NOR2XL inst_cellmath__24_0_I1045 (.Y(N4724), .A(N4395), .B(N4715));
NOR2XL inst_cellmath__24_0_I1046 (.Y(N3559), .A(N4395), .B(N4184));
NOR2XL inst_cellmath__24_0_I1047 (.Y(N4464), .A(N4395), .B(N3666));
NOR2XL inst_cellmath__24_0_I1048 (.Y(N3290), .A(N4395), .B(N3133));
NOR2XL inst_cellmath__24_0_I1049 (.Y(N4196), .A(N4395), .B(N4672));
NOR2XL inst_cellmath__24_0_I1050 (.Y(N5099), .A(N4395), .B(N4144));
INVXL inst_cellmath__24_0_I1051 (.Y(N3935), .A(N4395));
CLKINVX6 inst_cellmath__24_0_I1052 (.Y(N3861), .A(b_man[14]));
NOR2XL inst_cellmath__24_0_I1053 (.Y(N3595), .A(N3861), .B(N3346));
NOR2XL inst_cellmath__24_0_I1054 (.Y(N4497), .A(N3861), .B(N4891));
NOR2XL inst_cellmath__24_0_I1055 (.Y(N3322), .A(N3861), .B(N2934));
NOR2XL inst_cellmath__24_0_I1056 (.Y(N4231), .A(N3861), .B(N3835));
NOR2XL inst_cellmath__24_0_I1057 (.Y(N5131), .A(N3861), .B(N3299));
NOR2XL inst_cellmath__24_0_I1058 (.Y(N3967), .A(N4845), .B(N3861));
NOR2XL inst_cellmath__24_0_I1059 (.Y(N4871), .A(N3861), .B(N4318));
NOR2X1 inst_cellmath__24_0_I1060 (.Y(N3703), .A(N3861), .B(N3792));
NOR2X1 inst_cellmath__24_0_I1061 (.Y(N4604), .A(N3861), .B(N3260));
NOR2X1 inst_cellmath__24_0_I1062 (.Y(N3441), .A(N4801), .B(N3861));
NOR2X1 inst_cellmath__24_0_I1063 (.Y(N4338), .A(N3861), .B(N4273));
NOR2X1 inst_cellmath__24_0_I1064 (.Y(N3172), .A(N3751), .B(N3861));
NOR2XL inst_cellmath__24_0_I1065 (.Y(N4079), .A(N3861), .B(N3220));
NOR2X1 inst_cellmath__24_0_I1066 (.Y(N4982), .A(N3861), .B(N4758));
NOR2XL inst_cellmath__24_0_I1067 (.Y(N3814), .A(N3861), .B(N4232));
NOR2XL inst_cellmath__24_0_I1068 (.Y(N4714), .A(N3861), .B(N3704));
NOR2XL inst_cellmath__24_0_I1069 (.Y(N3549), .A(N3861), .B(N3176));
NOR2XL inst_cellmath__24_0_I1070 (.Y(N4453), .A(N3861), .B(N4715));
NOR2XL inst_cellmath__24_0_I1071 (.Y(N3282), .A(N3861), .B(N4184));
NOR2XL inst_cellmath__24_0_I1072 (.Y(N4183), .A(N3861), .B(N3666));
NOR2XL inst_cellmath__24_0_I1073 (.Y(N5089), .A(N3861), .B(N3133));
NOR2XL inst_cellmath__24_0_I1074 (.Y(N3926), .A(N3861), .B(N4672));
NOR2XL inst_cellmath__24_0_I1075 (.Y(N4824), .A(N3861), .B(N4144));
INVXL inst_cellmath__24_0_I1076 (.Y(N3662), .A(N3861));
CLKINVX6 inst_cellmath__24_0_I1077 (.Y(N4955), .A(b_man[15]));
NOR2XL inst_cellmath__24_0_I1078 (.Y(N3313), .A(N4955), .B(N3346));
NOR2XL inst_cellmath__24_0_I1079 (.Y(N4216), .A(N4955), .B(N4891));
NOR2XL inst_cellmath__24_0_I1080 (.Y(N5123), .A(N4955), .B(N2934));
NOR2XL inst_cellmath__24_0_I1081 (.Y(N3957), .A(N4955), .B(N3835));
NOR2X2 inst_cellmath__24_0_I1082 (.Y(N4858), .A(N3299), .B(N4955));
NOR2XL inst_cellmath__24_0_I1083 (.Y(N3694), .A(N4845), .B(N4955));
NOR2X1 inst_cellmath__24_0_I1084 (.Y(N4595), .A(N4955), .B(N4318));
NOR2X2 inst_cellmath__24_0_I1085 (.Y(N3430), .A(N3792), .B(N4955));
NOR2XL inst_cellmath__24_0_I1086 (.Y(N4330), .A(N4955), .B(N3260));
NOR2X1 inst_cellmath__24_0_I1087 (.Y(N3162), .A(N4801), .B(N4955));
NOR2X1 inst_cellmath__24_0_I1088 (.Y(N4069), .A(N4955), .B(N4273));
NOR2XL inst_cellmath__24_0_I1089 (.Y(N4973), .A(N4955), .B(N3751));
NOR2XL inst_cellmath__24_0_I1090 (.Y(N3805), .A(N4955), .B(N3220));
NOR2XL inst_cellmath__24_0_I1091 (.Y(N4705), .A(N4955), .B(N4758));
NOR2XL inst_cellmath__24_0_I1092 (.Y(N3541), .A(N4955), .B(N4232));
NOR2XL inst_cellmath__24_0_I1093 (.Y(N4445), .A(N4955), .B(N3704));
NOR2XL inst_cellmath__24_0_I1094 (.Y(N3273), .A(N4955), .B(N3176));
NOR2XL inst_cellmath__24_0_I1095 (.Y(N4175), .A(N4955), .B(N4715));
NOR2XL inst_cellmath__24_0_I1096 (.Y(N5081), .A(N4955), .B(N4184));
NOR2XL inst_cellmath__24_0_I1097 (.Y(N3915), .A(N4955), .B(N3666));
NOR2XL inst_cellmath__24_0_I1098 (.Y(N4814), .A(N4955), .B(N3133));
NOR2XL inst_cellmath__24_0_I1099 (.Y(N3651), .A(N4955), .B(N4672));
NOR2XL inst_cellmath__24_0_I1100 (.Y(N4557), .A(N4955), .B(N4144));
INVXL inst_cellmath__24_0_I1101 (.Y(N3387), .A(N4955));
CLKINVX12 inst_cellmath__24_0_I1102 (.Y(N3978), .A(b_man[16]));
NOR2XL inst_cellmath__24_0_I1103 (.Y(N5114), .A(N3978), .B(N3346));
NOR2XL inst_cellmath__24_0_I1104 (.Y(N3946), .A(N3978), .B(N4891));
NOR2XL inst_cellmath__24_0_I1105 (.Y(N4847), .A(N3978), .B(N2934));
NOR2X1 inst_cellmath__24_0_I1106 (.Y(N3687), .A(N3978), .B(N3835));
NOR2XL inst_cellmath__24_0_I1107 (.Y(N4586), .A(N3978), .B(N3299));
NOR2XL inst_cellmath__24_0_I1108 (.Y(N3419), .A(N3978), .B(N4845));
NOR2X2 inst_cellmath__24_0_I1109 (.Y(N4323), .A(N4318), .B(N3978));
NOR2X2 inst_cellmath__24_0_I1110 (.Y(N3154), .A(N3792), .B(N3978));
NOR2X1 inst_cellmath__24_0_I1111 (.Y(N4059), .A(N3978), .B(N3260));
NOR2X1 inst_cellmath__24_0_I1112 (.Y(N4964), .A(N3978), .B(N4801));
NOR2XL inst_cellmath__24_0_I1113 (.Y(N3797), .A(N3978), .B(N4273));
NOR2XL inst_cellmath__24_0_I1114 (.Y(N4695), .A(N3978), .B(N3751));
NOR2XL inst_cellmath__24_0_I1115 (.Y(N3536), .A(N3220), .B(N3978));
NOR2XL inst_cellmath__24_0_I1116 (.Y(N4436), .A(N3978), .B(N4758));
NOR2XL inst_cellmath__24_0_I1117 (.Y(N3263), .A(N3978), .B(N4232));
NOR2XL inst_cellmath__24_0_I1118 (.Y(N4169), .A(N3978), .B(N3704));
NOR2XL inst_cellmath__24_0_I1119 (.Y(N5071), .A(N3978), .B(N3176));
NOR2XL inst_cellmath__24_0_I1120 (.Y(N3905), .A(N3978), .B(N4715));
NOR2XL inst_cellmath__24_0_I1121 (.Y(N4805), .A(N3978), .B(N4184));
NOR2XL inst_cellmath__24_0_I1122 (.Y(N3641), .A(N3978), .B(N3666));
NOR2XL inst_cellmath__24_0_I1123 (.Y(N4549), .A(N3978), .B(N3133));
NOR2XL inst_cellmath__24_0_I1124 (.Y(N3375), .A(N3978), .B(N4672));
NOR2XL inst_cellmath__24_0_I1125 (.Y(N4278), .A(N3978), .B(N4144));
INVXL inst_cellmath__24_0_I1126 (.Y(N3116), .A(N3978));
CLKINVX12 inst_cellmath__24_0_I1127 (.Y(N3448), .A(b_man[17]));
NOR2XL inst_cellmath__24_0_I1128 (.Y(N4838), .A(N3448), .B(N3346));
NOR2XL inst_cellmath__24_0_I1129 (.Y(N3680), .A(N3448), .B(N4891));
NOR2XL inst_cellmath__24_0_I1130 (.Y(N4576), .A(N3448), .B(N2934));
NOR2XL inst_cellmath__24_0_I1131 (.Y(N3409), .A(N3448), .B(N3835));
NOR2X1 inst_cellmath__24_0_I1132 (.Y(N4315), .A(N3299), .B(N3448));
NOR2X1 inst_cellmath__24_0_I1133 (.Y(N3145), .A(N4845), .B(N3448));
NOR2X4 inst_cellmath__24_0_I1134 (.Y(N4051), .A(N3448), .B(N4318));
NOR2X2 inst_cellmath__24_0_I1135 (.Y(N4954), .A(N3448), .B(N3792));
NOR2X1 inst_cellmath__24_0_I1136 (.Y(N3789), .A(N3448), .B(N3260));
NOR2XL inst_cellmath__24_0_I1137 (.Y(N4685), .A(N3448), .B(N4801));
NOR2X1 inst_cellmath__24_0_I1138 (.Y(N3528), .A(N3448), .B(N4273));
NOR2XL inst_cellmath__24_0_I1139 (.Y(N4426), .A(N3448), .B(N3751));
NOR2XL inst_cellmath__24_0_I1140 (.Y(N3254), .A(N3448), .B(N3220));
NOR2XL inst_cellmath__24_0_I1141 (.Y(N4160), .A(N3448), .B(N4758));
NOR2XL inst_cellmath__24_0_I1142 (.Y(N5065), .A(N3448), .B(N4232));
NOR2XL inst_cellmath__24_0_I1143 (.Y(N3893), .A(N3448), .B(N3704));
NOR2XL inst_cellmath__24_0_I1144 (.Y(N4797), .A(N3448), .B(N3176));
NOR2XL inst_cellmath__24_0_I1145 (.Y(N3634), .A(N3448), .B(N4715));
NOR2XL inst_cellmath__24_0_I1146 (.Y(N4536), .A(N3448), .B(N4184));
NOR2XL inst_cellmath__24_0_I1147 (.Y(N3366), .A(N3448), .B(N3666));
NOR2XL inst_cellmath__24_0_I1148 (.Y(N4267), .A(N3448), .B(N3133));
NOR2XL inst_cellmath__24_0_I1149 (.Y(N3103), .A(N3448), .B(N4672));
NOR2XL inst_cellmath__24_0_I1150 (.Y(N4012), .A(N3448), .B(N4144));
INVXL inst_cellmath__24_0_I1151 (.Y(N4909), .A(N3448));
CLKINVX8 inst_cellmath__24_0_I1152 (.Y(N4990), .A(b_man[18]));
NOR2XL inst_cellmath__24_0_I1154 (.Y(N4569), .A(N4990), .B(N3346));
NOR2XL inst_cellmath__24_0_I1155 (.Y(N3399), .A(N4891), .B(N4990));
NOR2XL inst_cellmath__24_0_I1156 (.Y(N4305), .A(N4990), .B(N2934));
NOR2X1 inst_cellmath__24_0_I1157 (.Y(N3137), .A(N4990), .B(N3835));
NOR2X2 inst_cellmath__24_0_I1158 (.Y(N4042), .A(N3299), .B(N4990));
NOR2X1 inst_cellmath__24_0_I1159 (.Y(N4945), .A(N4845), .B(N4990));
NOR2X2 inst_cellmath__24_0_I1160 (.Y(N3780), .A(N4990), .B(N4318));
NOR2XL inst_cellmath__24_0_I1161 (.Y(N4676), .A(N4990), .B(N3792));
NOR2XL inst_cellmath__24_0_I1162 (.Y(N3519), .A(N4990), .B(N3260));
NOR2XL inst_cellmath__24_0_I1163 (.Y(N4417), .A(N4990), .B(N4801));
NOR2X1 inst_cellmath__24_0_I1164 (.Y(N3245), .A(N4990), .B(N4273));
NOR2XL inst_cellmath__24_0_I1165 (.Y(N4150), .A(N3751), .B(N4990));
NOR2XL inst_cellmath__24_0_I1166 (.Y(N5055), .A(N4990), .B(N3220));
NOR2XL inst_cellmath__24_0_I1167 (.Y(N3885), .A(N4990), .B(N4758));
NOR2XL inst_cellmath__24_0_I1168 (.Y(N4787), .A(N4990), .B(N4232));
NOR2XL inst_cellmath__24_0_I1169 (.Y(N3626), .A(N4990), .B(N3704));
NOR2XL inst_cellmath__24_0_I1170 (.Y(N4526), .A(N4990), .B(N3176));
NOR2XL inst_cellmath__24_0_I1171 (.Y(N3356), .A(N4990), .B(N4715));
NOR2XL inst_cellmath__24_0_I1172 (.Y(N4258), .A(N4990), .B(N4184));
NOR2XL inst_cellmath__24_0_I1173 (.Y(N3094), .A(N4990), .B(N3666));
NOR2XL inst_cellmath__24_0_I1174 (.Y(N4001), .A(N4990), .B(N3133));
NOR2XL inst_cellmath__24_0_I1175 (.Y(N4901), .A(N4990), .B(N4672));
NOR2XL inst_cellmath__24_0_I1176 (.Y(N3735), .A(N4990), .B(N4144));
INVXL inst_cellmath__24_0_I1177 (.Y(N4635), .A(N4990));
CLKINVX6 inst_cellmath__24_0_I1178 (.Y(N4463), .A(b_man[19]));
NOR2XL inst_cellmath__24_0_I1179 (.Y(N4295), .A(N4463), .B(N3346));
NOR2XL inst_cellmath__24_0_I1180 (.Y(N3129), .A(N4463), .B(N4891));
NOR2XL inst_cellmath__24_0_I1181 (.Y(N4035), .A(N4463), .B(N2934));
NOR2X2 inst_cellmath__24_0_I1182 (.Y(N4938), .A(N3835), .B(N4463));
NOR2X2 inst_cellmath__24_0_I1183 (.Y(N3773), .A(N3299), .B(N4463));
NOR2X1 inst_cellmath__24_0_I1184 (.Y(N4667), .A(N4463), .B(N4845));
NOR2X1 inst_cellmath__24_0_I5206 (.Y(N11813), .A(N4463), .B(N4318));
NOR2XL inst_cellmath__24_0_I1186 (.Y(N4409), .A(N4463), .B(N3792));
NOR2XL inst_cellmath__24_0_I1187 (.Y(N3238), .A(N4463), .B(N3260));
NOR2XL inst_cellmath__24_0_I1188 (.Y(N4141), .A(N4463), .B(N4801));
NOR2XL inst_cellmath__24_0_I1189 (.Y(N5047), .A(N4463), .B(N4273));
NOR2XL inst_cellmath__24_0_I1190 (.Y(N3876), .A(N4463), .B(N3751));
NOR2XL inst_cellmath__24_0_I1191 (.Y(N4779), .A(N4463), .B(N3220));
NOR2XL inst_cellmath__24_0_I1192 (.Y(N3617), .A(N4463), .B(N4758));
NOR2XL inst_cellmath__24_0_I1193 (.Y(N4518), .A(N4463), .B(N4232));
NOR2XL inst_cellmath__24_0_I1194 (.Y(N3348), .A(N4463), .B(N3704));
NOR2XL inst_cellmath__24_0_I1195 (.Y(N4250), .A(N4463), .B(N3176));
NOR2XL inst_cellmath__24_0_I1196 (.Y(N3085), .A(N4463), .B(N4715));
NOR2XL inst_cellmath__24_0_I1197 (.Y(N3992), .A(N4463), .B(N4184));
NOR2XL inst_cellmath__24_0_I1198 (.Y(N4893), .A(N4463), .B(N3666));
NOR2XL inst_cellmath__24_0_I1199 (.Y(N3727), .A(N4463), .B(N3133));
NOR2XL inst_cellmath__24_0_I1200 (.Y(N4626), .A(N4463), .B(N4672));
NOR2XL inst_cellmath__24_0_I1201 (.Y(N3464), .A(N4463), .B(N4144));
INVXL inst_cellmath__24_0_I1202 (.Y(N4362), .A(N4463));
CLKINVX6 inst_cellmath__24_0_I1203 (.Y(N3931), .A(b_man[20]));
NOR2XL inst_cellmath__24_0_I1204 (.Y(N4025), .A(N3931), .B(N3346));
NOR2XL inst_cellmath__24_0_I1205 (.Y(N4926), .A(N3931), .B(N4891));
NOR2XL inst_cellmath__24_0_I1206 (.Y(N3762), .A(N3931), .B(N2934));
NOR2X4 inst_cellmath__24_0_I1207 (.Y(N4659), .A(N3931), .B(N3835));
NOR2X1 inst_cellmath__24_0_I1208 (.Y(N3500), .A(N3299), .B(N3931));
NOR2X1 inst_cellmath__24_0_I1209 (.Y(N4402), .A(N4845), .B(N3931));
NOR2XL inst_cellmath__24_0_I1210 (.Y(N3230), .A(N3931), .B(N4318));
NOR2XL inst_cellmath__24_0_I1211 (.Y(N4133), .A(N3931), .B(N3792));
NOR2XL inst_cellmath__24_0_I1212 (.Y(N5039), .A(N3931), .B(N3260));
NOR2XL inst_cellmath__24_0_I1213 (.Y(N3869), .A(N3931), .B(N4801));
NOR2XL inst_cellmath__24_0_I1214 (.Y(N4770), .A(N3931), .B(N4273));
NOR2XL inst_cellmath__24_0_I1215 (.Y(N3608), .A(N3931), .B(N3751));
NOR2XL inst_cellmath__24_0_I1216 (.Y(N4508), .A(N3931), .B(N3220));
NOR2XL inst_cellmath__24_0_I1217 (.Y(N3340), .A(N3931), .B(N4758));
NOR2XL inst_cellmath__24_0_I1218 (.Y(N4243), .A(N3931), .B(N4232));
NOR2XL inst_cellmath__24_0_I1219 (.Y(N5144), .A(N3931), .B(N3704));
NOR2XL inst_cellmath__24_0_I1220 (.Y(N3983), .A(N3931), .B(N3176));
NOR2XL inst_cellmath__24_0_I1221 (.Y(N4883), .A(N3931), .B(N4715));
NOR2XL inst_cellmath__24_0_I1222 (.Y(N3716), .A(N3931), .B(N4184));
NOR2XL inst_cellmath__24_0_I1223 (.Y(N4618), .A(N3931), .B(N3666));
NOR2XL inst_cellmath__24_0_I1224 (.Y(N3453), .A(N3931), .B(N3133));
NOR2XL inst_cellmath__24_0_I1225 (.Y(N4351), .A(N3931), .B(N4672));
NOR2XL inst_cellmath__24_0_I1226 (.Y(N3187), .A(N3931), .B(N4144));
INVXL inst_cellmath__24_0_I1227 (.Y(N4090), .A(N3931));
CLKINVX6 inst_cellmath__24_0_I1228 (.Y(N3404), .A(b_man[21]));
NOR2XL inst_cellmath__24_0_I1229 (.Y(N3754), .A(N3404), .B(N3346));
NOR2XL inst_cellmath__24_0_I1230 (.Y(N4649), .A(N3404), .B(N4891));
NOR2X1 inst_cellmath__24_0_I1231 (.Y(N3489), .A(N2934), .B(N3404));
NOR2X1 inst_cellmath__24_0_I1232 (.Y(N4391), .A(N3404), .B(N3835));
NOR2XL inst_cellmath__24_0_I1233 (.Y(N3222), .A(N3404), .B(N3299));
NOR2XL inst_cellmath__24_0_I1234 (.Y(N4124), .A(N3404), .B(N4845));
NOR2XL inst_cellmath__24_0_I1235 (.Y(N5031), .A(N3404), .B(N4318));
NOR2XL inst_cellmath__24_0_I1236 (.Y(N3859), .A(N3404), .B(N3792));
NOR2X1 inst_cellmath__24_0_I1237 (.Y(N4760), .A(N3404), .B(N3260));
NOR2XL inst_cellmath__24_0_I1238 (.Y(N3597), .A(N3404), .B(N4801));
NOR2XL inst_cellmath__24_0_I1239 (.Y(N4501), .A(N3404), .B(N4273));
NOR2XL inst_cellmath__24_0_I1240 (.Y(N3326), .A(N3404), .B(N3751));
NOR2XL inst_cellmath__24_0_I1241 (.Y(N4234), .A(N3404), .B(N3220));
NOR2XL inst_cellmath__24_0_I1242 (.Y(N5135), .A(N3404), .B(N4758));
NOR2XL inst_cellmath__24_0_I1243 (.Y(N3971), .A(N3404), .B(N4232));
NOR2XL inst_cellmath__24_0_I1244 (.Y(N4873), .A(N3404), .B(N3704));
NOR2XL inst_cellmath__24_0_I1245 (.Y(N3707), .A(N3404), .B(N3176));
NOR2XL inst_cellmath__24_0_I1246 (.Y(N4607), .A(N3404), .B(N4715));
NOR2XL inst_cellmath__24_0_I1247 (.Y(N3443), .A(N3404), .B(N4184));
NOR2XL inst_cellmath__24_0_I1248 (.Y(N4340), .A(N3404), .B(N3666));
NOR2XL inst_cellmath__24_0_I1249 (.Y(N3178), .A(N3404), .B(N3133));
NOR2XL inst_cellmath__24_0_I1250 (.Y(N4081), .A(N3404), .B(N4672));
NOR2XL inst_cellmath__24_0_I1251 (.Y(N4984), .A(N3404), .B(N4144));
INVXL inst_cellmath__24_0_I1252 (.Y(N3818), .A(N3404));
INVX3 inst_cellmath__24_0_I1253 (.Y(N4946), .A(b_man[22]));
NOR2XL inst_cellmath__24_0_I1254 (.Y(N3477), .A(N4946), .B(N3346));
NOR2XL inst_cellmath__24_0_I1255 (.Y(N4380), .A(N4946), .B(N4891));
NOR2XL inst_cellmath__24_0_I1256 (.Y(N3211), .A(N4946), .B(N2934));
NOR2XL inst_cellmath__24_0_I1257 (.Y(N4113), .A(N4946), .B(N3835));
NOR2XL inst_cellmath__24_0_I1258 (.Y(N5021), .A(N4946), .B(N3299));
NOR2XL inst_cellmath__24_0_I1259 (.Y(N3851), .A(N4946), .B(N4845));
NOR2XL inst_cellmath__24_0_I1260 (.Y(N4750), .A(N4946), .B(N4318));
NOR2XL inst_cellmath__24_0_I1261 (.Y(N3587), .A(N4946), .B(N3792));
NOR2XL inst_cellmath__24_0_I1262 (.Y(N4493), .A(N4946), .B(N3260));
NOR2XL inst_cellmath__24_0_I1263 (.Y(N3317), .A(N4946), .B(N4801));
NOR2XL inst_cellmath__24_0_I1264 (.Y(N4222), .A(N4946), .B(N4273));
NOR2XL inst_cellmath__24_0_I1265 (.Y(N5125), .A(N4946), .B(N3751));
NOR2XL inst_cellmath__24_0_I1266 (.Y(N3961), .A(N4946), .B(N3220));
NOR2XL inst_cellmath__24_0_I1267 (.Y(N4864), .A(N4946), .B(N4758));
NOR2XL inst_cellmath__24_0_I1268 (.Y(N3697), .A(N4946), .B(N4232));
NOR2XL inst_cellmath__24_0_I1269 (.Y(N4598), .A(N4946), .B(N3704));
NOR2XL inst_cellmath__24_0_I1270 (.Y(N3433), .A(N4946), .B(N3176));
NOR2XL inst_cellmath__24_0_I1271 (.Y(N4332), .A(N4946), .B(N4715));
NOR2XL inst_cellmath__24_0_I1272 (.Y(N3165), .A(N4946), .B(N4184));
NOR2XL inst_cellmath__24_0_I1273 (.Y(N4072), .A(N4946), .B(N3666));
NOR2XL inst_cellmath__24_0_I1274 (.Y(N4977), .A(N4946), .B(N3133));
NOR2XL inst_cellmath__24_0_I1275 (.Y(N3808), .A(N4946), .B(N4672));
NOR2XL inst_cellmath__24_0_I1276 (.Y(N4708), .A(N4946), .B(N4144));
INVXL inst_cellmath__24_0_I1277 (.Y(N3544), .A(N4946));
INVXL inst_cellmath__24_0_I1278 (.Y(N3468), .A(N3346));
INVX1 inst_cellmath__24_0_I1279 (.Y(N4371), .A(N4891));
INVX1 inst_cellmath__24_0_I1280 (.Y(N3201), .A(N2934));
INVXL inst_cellmath__24_0_I1281 (.Y(N4104), .A(N3835));
INVXL inst_cellmath__24_0_I1282 (.Y(N5012), .A(N3299));
INVXL inst_cellmath__24_0_I1283 (.Y(N3842), .A(N4845));
INVXL inst_cellmath__24_0_I1284 (.Y(N4740), .A(N4318));
INVXL inst_cellmath__24_0_I1285 (.Y(N3579), .A(N3792));
INVXL inst_cellmath__24_0_I1286 (.Y(N4483), .A(N3260));
INVXL inst_cellmath__24_0_I1287 (.Y(N3307), .A(N4801));
INVXL inst_cellmath__24_0_I1288 (.Y(N4213), .A(N4273));
INVXL inst_cellmath__24_0_I1289 (.Y(N5116), .A(N3751));
INVXL inst_cellmath__24_0_I1290 (.Y(N3951), .A(N3220));
INVXL inst_cellmath__24_0_I1291 (.Y(N4854), .A(N4758));
INVXL inst_cellmath__24_0_I1292 (.Y(N3689), .A(N4232));
INVXL inst_cellmath__24_0_I1293 (.Y(N4590), .A(N3704));
INVXL inst_cellmath__24_0_I1294 (.Y(N3425), .A(N3176));
INVXL inst_cellmath__24_0_I1295 (.Y(N4326), .A(N4715));
INVXL inst_cellmath__24_0_I1296 (.Y(N3157), .A(N4184));
INVXL inst_cellmath__24_0_I1297 (.Y(N4063), .A(N3666));
INVXL inst_cellmath__24_0_I1298 (.Y(N4967), .A(N3133));
INVXL inst_cellmath__24_0_I1299 (.Y(N3801), .A(N4672));
INVXL inst_cellmath__24_0_I1300 (.Y(N4700), .A(N4144));
ADDHX1 inst_cellmath__24_0_I1301 (.CO(N4889), .S(N4440), .A(N5084), .B(N3907));
ADDHX1 inst_cellmath__24_0_I1302 (.CO(N3723), .S(N3268), .A(N3917), .B(N4807));
ADDFX1 inst_cellmath__24_0_I1303 (.CO(N4624), .S(N4171), .A(N4531), .B(N3637), .CI(N4889));
ADDHX1 inst_cellmath__24_0_I1304 (.CO(N3460), .S(N5076), .A(N4817), .B(N3646));
ADDFXL inst_cellmath__24_0_I1305 (.CO(N4358), .S(N3910), .A(N3358), .B(N4541), .CI(N4252));
ADDFXL inst_cellmath__24_0_I1306 (.CO(N3194), .S(N4809), .A(N3723), .B(N5076), .CI(N3910));
ADDHX1 inst_cellmath__24_0_I1307 (.CO(N4097), .S(N3645), .A(N3656), .B(N4550));
ADDFX1 inst_cellmath__24_0_I1308 (.CO(N5000), .S(N4552), .A(N4260), .B(N3367), .CI(N3087));
ADDFX1 inst_cellmath__24_0_I1309 (.CO(N3834), .S(N3380), .A(N3460), .B(N3985), .CI(N3645));
ADDFX1 inst_cellmath__24_0_I1310 (.CO(N4730), .S(N4282), .A(N4552), .B(N4358), .CI(N3194));
ADDHX1 inst_cellmath__24_0_I1311 (.CO(N3568), .S(N3119), .A(N4558), .B(N3378));
ADDFXL inst_cellmath__24_0_I1312 (.CO(N4475), .S(N4021), .A(N3097), .B(N4272), .CI(N3993));
ADDFX1 inst_cellmath__24_0_I1313 (.CO(N3297), .S(N4925), .A(N3711), .B(N4886), .CI(N4097));
ADDFXL inst_cellmath__24_0_I1314 (.CO(N4206), .S(N3759), .A(N5000), .B(N3119), .CI(N4021));
ADDFX1 inst_cellmath__24_0_I1315 (.CO(N5108), .S(N4654), .A(N4925), .B(N3834), .CI(N3759));
ADDHX1 inst_cellmath__24_0_I1316 (.CO(N3941), .S(N3499), .A(N3389), .B(N4283));
ADDFX1 inst_cellmath__24_0_I1317 (.CO(N4844), .S(N4398), .A(N4003), .B(N3108), .CI(N4895));
ADDFX1 inst_cellmath__24_0_I1318 (.CO(N3682), .S(N3226), .A(N4609), .B(N3720), .CI(N3435));
ADDFX1 inst_cellmath__24_0_I1319 (.CO(N4579), .S(N4132), .A(N3499), .B(N3568), .CI(N4475));
ADDFX1 inst_cellmath__24_0_I1320 (.CO(N3416), .S(N5037), .A(N3226), .B(N4398), .CI(N3297));
ADDFX1 inst_cellmath__24_0_I1321 (.CO(N4317), .S(N3863), .A(N4132), .B(N4206), .CI(N5037));
ADDHXL inst_cellmath__24_0_I1322 (.CO(N3148), .S(N4768), .A(N4292), .B(N3117));
ADDFXL inst_cellmath__24_0_I1323 (.CO(N4057), .S(N3603), .A(N4903), .B(N4013), .CI(N3729));
ADDFXL inst_cellmath__24_0_I1324 (.CO(N4957), .S(N4504), .A(N4335), .B(N4619), .CI(N3444));
ADDFXL inst_cellmath__24_0_I1325 (.CO(N3791), .S(N3338), .A(N3160), .B(N3941), .CI(N4768));
ADDFX1 inst_cellmath__24_0_I1326 (.CO(N4691), .S(N4240), .A(N3682), .B(N4844), .CI(N3603));
ADDFX1 inst_cellmath__24_0_I1327 (.CO(N3530), .S(N5140), .A(N4579), .B(N4504), .CI(N3338));
ADDFX1 inst_cellmath__24_0_I1328 (.CO(N4428), .S(N3981), .A(N4240), .B(N3416), .CI(N5140));
ADDHX1 inst_cellmath__24_0_I1329 (.CO(N3259), .S(N4879), .A(N3124), .B(N4022));
ADDFX1 inst_cellmath__24_0_I1330 (.CO(N4162), .S(N3713), .A(N3738), .B(N4914), .CI(N4627));
ADDFX1 inst_cellmath__24_0_I1331 (.CO(N5067), .S(N4616), .A(N4345), .B(N3458), .CI(N3168));
ADDFX1 inst_cellmath__24_0_I1332 (.CO(N3899), .S(N3450), .A(N4960), .B(N4064), .CI(N3148));
ADDFXL inst_cellmath__24_0_I1333 (.CO(N4800), .S(N4347), .A(N4879), .B(N4957), .CI(N4057));
ADDFX1 inst_cellmath__24_0_I1334 (.CO(N3636), .S(N3185), .A(N4616), .B(N3713), .CI(N3791));
ADDFXL inst_cellmath__24_0_I1335 (.CO(N4544), .S(N4087), .A(N4691), .B(N3450), .CI(N4347));
ADDFXL inst_cellmath__24_0_I1336 (.CO(N3369), .S(N4992), .A(N3185), .B(N3530), .CI(N4087));
ADDHX1 inst_cellmath__24_0_I1337 (.CO(N4271), .S(N3826), .A(N4031), .B(N4923));
ADDFX1 inst_cellmath__24_0_I1338 (.CO(N3111), .S(N4723), .A(N4636), .B(N3748), .CI(N3466));
ADDFX1 inst_cellmath__24_0_I1339 (.CO(N4015), .S(N3558), .A(N3179), .B(N4354), .CI(N4073));
ADDFX1 inst_cellmath__24_0_I1340 (.CO(N4913), .S(N4466), .A(N3794), .B(N4970), .CI(N4683));
ADDFX1 inst_cellmath__24_0_I1341 (.CO(N3750), .S(N3289), .A(N3826), .B(N3259), .CI(N4162));
ADDFHXL inst_cellmath__24_0_I1342 (.CO(N4647), .S(N4195), .A(N5067), .B(N3899), .CI(N4723));
ADDFX1 inst_cellmath__24_0_I1343 (.CO(N3485), .S(N5101), .A(N4466), .B(N3558), .CI(N4800));
ADDFX1 inst_cellmath__24_0_I1344 (.CO(N4387), .S(N3934), .A(N3636), .B(N3289), .CI(N4195));
ADDFHXL inst_cellmath__24_0_I1345 (.CO(N3218), .S(N4834), .A(N4544), .B(N5101), .CI(N3934));
ADDHX1 inst_cellmath__24_0_I1346 (.CO(N4121), .S(N3674), .A(N3757), .B(N4932));
ADDFX1 inst_cellmath__24_0_I1347 (.CO(N5028), .S(N4573), .A(N4645), .B(N3475), .CI(N4365));
ADDFX1 inst_cellmath__24_0_I1348 (.CO(N3856), .S(N3405), .A(N4082), .B(N3188), .CI(N4980));
ADDFX1 inst_cellmath__24_0_I1349 (.CO(N4756), .S(N4308), .A(N4692), .B(N3803), .CI(N3523));
ADDFX1 inst_cellmath__24_0_I1350 (.CO(N3594), .S(N3141), .A(N4271), .B(N4414), .CI(N3674));
ADDFXL inst_cellmath__24_0_I1351 (.CO(N4496), .S(N4048), .A(N4913), .B(N4015), .CI(N3111));
ADDFXL inst_cellmath__24_0_I1352 (.CO(N3325), .S(N4949), .A(N4308), .B(N3405), .CI(N4573));
ADDFX1 inst_cellmath__24_0_I1353 (.CO(N4230), .S(N3783), .A(N3141), .B(N3750), .CI(N4048));
ADDFXL inst_cellmath__24_0_I1354 (.CO(N5130), .S(N4682), .A(N3485), .B(N4647), .CI(N4949));
ADDFXL inst_cellmath__24_0_I1355 (.CO(N3970), .S(N3522), .A(N3783), .B(N4387), .CI(N4682));
ADDHX1 inst_cellmath__24_0_I1356 (.CO(N4870), .S(N4419), .A(N3767), .B(N4655));
ADDFXL inst_cellmath__24_0_I1357 (.CO(N3702), .S(N3251), .A(N4374), .B(N3486), .CI(N3196));
ADDFX1 inst_cellmath__24_0_I1358 (.CO(N4606), .S(N4154), .A(N4989), .B(N4094), .CI(N3811));
ADDFX1 inst_cellmath__24_0_I1359 (.CO(N3440), .S(N5057), .A(N3533), .B(N4701), .CI(N4422));
ADDFX1 inst_cellmath__24_0_I1360 (.CO(N4337), .S(N3890), .A(N4137), .B(N3242), .CI(N4121));
ADDFX1 inst_cellmath__24_0_I1361 (.CO(N3175), .S(N4790), .A(N5028), .B(N4419), .CI(N3856));
ADDFX1 inst_cellmath__24_0_I1362 (.CO(N4078), .S(N3627), .A(N4756), .B(N3251), .CI(N4154));
ADDFX1 inst_cellmath__24_0_I1363 (.CO(N4981), .S(N4533), .A(N3594), .B(N5057), .CI(N4496));
ADDFX1 inst_cellmath__24_0_I1364 (.CO(N3816), .S(N3360), .A(N3325), .B(N3890), .CI(N4790));
ADDFX1 inst_cellmath__24_0_I1365 (.CO(N4713), .S(N4259), .A(N4533), .B(N3627), .CI(N4230));
ADDFX1 inst_cellmath__24_0_I1366 (.CO(N3548), .S(N3099), .A(N5130), .B(N3360), .CI(N4259));
ADDHX1 inst_cellmath__24_0_I1367 (.CO(N4456), .S(N4005), .A(N4664), .B(N3496));
ADDFXL inst_cellmath__24_0_I1368 (.CO(N3281), .S(N4902), .A(N3206), .B(N4385), .CI(N4102));
ADDFX1 inst_cellmath__24_0_I1369 (.CO(N4182), .S(N3741), .A(N3819), .B(N11781), .CI(N4709));
ADDFX1 inst_cellmath__24_0_I1370 (.CO(N5091), .S(N4638), .A(N3539), .B(N3252), .CI(N4432));
ADDFX1 inst_cellmath__24_0_I1371 (.CO(N3925), .S(N3474), .A(N5044), .B(N4145), .CI(N3864));
ADDFX1 inst_cellmath__24_0_I1372 (.CO(N4823), .S(N4377), .A(N4005), .B(N4870), .CI(N3702));
ADDFX1 inst_cellmath__24_0_I1373 (.CO(N3665), .S(N3208), .A(N3440), .B(N4606), .CI(N4902));
ADDFXL inst_cellmath__24_0_I1374 (.CO(N4565), .S(N4110), .A(N4638), .B(N4337), .CI(N3741));
ADDFXL inst_cellmath__24_0_I1375 (.CO(N3396), .S(N5018), .A(N3175), .B(N3474), .CI(N4078));
ADDFX1 inst_cellmath__24_0_I1376 (.CO(N4300), .S(N3849), .A(N4377), .B(N3208), .CI(N4110));
ADDFXL inst_cellmath__24_0_I1377 (.CO(N3132), .S(N4747), .A(N3816), .B(N4981), .CI(N5018));
ADDFXL inst_cellmath__24_0_I1378 (.CO(N4038), .S(N3585), .A(N4713), .B(N3849), .CI(N4747));
ADDHXL inst_cellmath__24_0_I1379 (.CO(N4940), .S(N4490), .A(N3505), .B(N4396));
ADDFX1 inst_cellmath__24_0_I1380 (.CO(N3776), .S(N3312), .A(N3216), .B(N4111), .CI(N5005));
ADDFX1 inst_cellmath__24_0_I1381 (.CO(N4671), .S(N4220), .A(N4718), .B(N3829), .CI(N3547));
ADDFX1 inst_cellmath__24_0_I1382 (.CO(N3513), .S(N5122), .A(N3261), .B(N4443), .CI(N4156));
ADDFX1 inst_cellmath__24_0_I1383 (.CO(N4411), .S(N3956), .A(N3873), .B(N5052), .CI(N4765));
ADDFX1 inst_cellmath__24_0_I1384 (.CO(N3240), .S(N4861), .A(N4456), .B(N3595), .CI(N4490));
ADDFXL inst_cellmath__24_0_I1385 (.CO(N4143), .S(N3693), .A(N5091), .B(N4182), .CI(N3281));
ADDFX1 inst_cellmath__24_0_I1386 (.CO(N5050), .S(N4594), .A(N3312), .B(N3925), .CI(N4220));
ADDFX1 inst_cellmath__24_0_I1387 (.CO(N3878), .S(N3429), .A(N3956), .B(N5122), .CI(N4823));
ADDFX1 inst_cellmath__24_0_I1388 (.CO(N4781), .S(N4329), .A(N4861), .B(N3665), .CI(N3693));
ADDFX1 inst_cellmath__24_0_I1389 (.CO(N3619), .S(N3164), .A(N4594), .B(N4565), .CI(N3396));
ADDFHXL inst_cellmath__24_0_I1390 (.CO(N4521), .S(N4068), .A(N3429), .B(N4300), .CI(N4329));
ADDFHXL inst_cellmath__24_0_I1391 (.CO(N3351), .S(N4972), .A(N3164), .B(N3132), .CI(N4068));
ADDHX1 inst_cellmath__24_0_I1392 (.CO(N4251), .S(N3807), .A(N4405), .B(N3227));
ADDFXL inst_cellmath__24_0_I1393 (.CO(N3089), .S(N4704), .A(N5016), .B(N4122), .CI(N3838));
ADDFX1 inst_cellmath__24_0_I1394 (.CO(N3995), .S(N3540), .A(N4451), .B(N4727), .CI(N3554));
ADDFX1 inst_cellmath__24_0_I1395 (.CO(N4894), .S(N4447), .A(N4165), .B(N3269), .CI(N5061));
ADDFX1 inst_cellmath__24_0_I1396 (.CO(N3731), .S(N3272), .A(N4774), .B(N3882), .CI(N3604));
ADDFX1 inst_cellmath__24_0_I1397 (.CO(N4629), .S(N4174), .A(N3313), .B(N4497), .CI(N4940));
ADDFX1 inst_cellmath__24_0_I1398 (.CO(N3465), .S(N5083), .A(N3807), .B(N3776), .CI(N4671));
ADDFXL inst_cellmath__24_0_I1399 (.CO(N4367), .S(N3914), .A(N4411), .B(N3513), .CI(N4704));
ADDFX1 inst_cellmath__24_0_I1400 (.CO(N3198), .S(N4813), .A(N4447), .B(N3540), .CI(N3272));
ADDFX1 inst_cellmath__24_0_I1401 (.CO(N4101), .S(N3654), .A(N4174), .B(N3240), .CI(N4143));
ADDFX1 inst_cellmath__24_0_I1402 (.CO(N5007), .S(N4556), .A(N5050), .B(N5083), .CI(N3914));
ADDFX1 inst_cellmath__24_0_I1403 (.CO(N3840), .S(N3386), .A(N3878), .B(N4813), .CI(N3654));
ADDFX1 inst_cellmath__24_0_I1404 (.CO(N4734), .S(N4290), .A(N4556), .B(N4781), .CI(N3619));
ADDFX1 inst_cellmath__24_0_I1405 (.CO(N3575), .S(N3123), .A(N4521), .B(N3386), .CI(N4290));
ADDHX1 inst_cellmath__24_0_I1406 (.CO(N4481), .S(N4028), .A(N3235), .B(N4130));
ADDFXL inst_cellmath__24_0_I1407 (.CO(N3302), .S(N4930), .A(N3847), .B(N5026), .CI(N4736));
ADDFX1 inst_cellmath__24_0_I1408 (.CO(N4210), .S(N3765), .A(N4458), .B(N3563), .CI(N3277));
ADDFX1 inst_cellmath__24_0_I1409 (.CO(N5113), .S(N4661), .A(N5069), .B(N4173), .CI(N3891));
ADDFX1 inst_cellmath__24_0_I1410 (.CO(N3945), .S(N3504), .A(N3614), .B(N4782), .CI(N4505));
ADDFX1 inst_cellmath__24_0_I1411 (.CO(N4850), .S(N4404), .A(N4216), .B(N3322), .CI(N5114));
ADDFX1 inst_cellmath__24_0_I1412 (.CO(N3686), .S(N3232), .A(N4028), .B(N4251), .CI(N3089));
ADDFX1 inst_cellmath__24_0_I1413 (.CO(N4585), .S(N4136), .A(N4894), .B(N3995), .CI(N3731));
ADDFXL inst_cellmath__24_0_I1414 (.CO(N3422), .S(N5041), .A(N4629), .B(N4930), .CI(N3765));
ADDFX1 inst_cellmath__24_0_I1415 (.CO(N4322), .S(N3870), .A(N3504), .B(N4661), .CI(N4404));
ADDFX1 inst_cellmath__24_0_I1416 (.CO(N3153), .S(N4773), .A(N4367), .B(N3465), .CI(N3198));
ADDFX1 inst_cellmath__24_0_I1417 (.CO(N4061), .S(N3611), .A(N3232), .B(N4136), .CI(N5041));
ADDFX1 inst_cellmath__24_0_I1418 (.CO(N4963), .S(N4511), .A(N4101), .B(N3870), .CI(N5007));
ADDFXL inst_cellmath__24_0_I1419 (.CO(N3796), .S(N3342), .A(N3611), .B(N4773), .CI(N3840));
ADDFX1 inst_cellmath__24_0_I1420 (.CO(N4697), .S(N4246), .A(N4734), .B(N4511), .CI(N3342));
ADDHXL inst_cellmath__24_0_I1421 (.CO(N3535), .S(N3079), .A(N4138), .B(N5035));
ADDFXL inst_cellmath__24_0_I1422 (.CO(N4435), .S(N3987), .A(N4748), .B(N3857), .CI(N3573));
ADDFX1 inst_cellmath__24_0_I1423 (.CO(N3265), .S(N4885), .A(N3287), .B(N4468), .CI(N4181));
ADDFX1 inst_cellmath__24_0_I1424 (.CO(N4168), .S(N3719), .A(N5079), .B(N4793), .CI(N3900));
ADDFXL inst_cellmath__24_0_I1425 (.CO(N5075), .S(N4621), .A(N4514), .B(N3623), .CI(N3334));
ADDFX1 inst_cellmath__24_0_I1426 (.CO(N3904), .S(N3457), .A(N5123), .B(N4231), .CI(N3946));
ADDFX1 inst_cellmath__24_0_I1427 (.CO(N4804), .S(N4357), .A(N4838), .B(N4481), .CI(N3079));
ADDFX1 inst_cellmath__24_0_I1428 (.CO(N3644), .S(N3190), .A(N5113), .B(N3302), .CI(N4210));
ADDFXL inst_cellmath__24_0_I1429 (.CO(N4548), .S(N4093), .A(N3945), .B(N4850), .CI(N3987));
ADDFXL inst_cellmath__24_0_I1430 (.CO(N3374), .S(N4999), .A(N3719), .B(N4621), .CI(N4885));
ADDFX1 inst_cellmath__24_0_I1431 (.CO(N4281), .S(N3831), .A(N4585), .B(N3457), .CI(N3686));
ADDFX1 inst_cellmath__24_0_I1432 (.CO(N3115), .S(N4726), .A(N3422), .B(N4357), .CI(N3190));
ADDFXL inst_cellmath__24_0_I1433 (.CO(N4018), .S(N3566), .A(N4322), .B(N4093), .CI(N4999));
ADDFXL inst_cellmath__24_0_I1434 (.CO(N4921), .S(N4470), .A(N3831), .B(N3153), .CI(N4061));
ADDFXL inst_cellmath__24_0_I1435 (.CO(N3756), .S(N3293), .A(N3566), .B(N4726), .CI(N4963));
ADDFXL inst_cellmath__24_0_I1436 (.CO(N4652), .S(N4202), .A(N3796), .B(N4470), .CI(N3293));
ADDHX1 inst_cellmath__24_0_I1437 (.CO(N3494), .S(N5106), .A(N5042), .B(N3865));
ADDFXL inst_cellmath__24_0_I1438 (.CO(N4394), .S(N3937), .A(N3582), .B(N4757), .CI(N4479));
ADDFX1 inst_cellmath__24_0_I1439 (.CO(N3224), .S(N4842), .A(N4190), .B(N5087), .CI(N3294));
ADDFX1 inst_cellmath__24_0_I1440 (.CO(N4129), .S(N3679), .A(N3629), .B(N3911), .CI(N4803));
ADDFX1 inst_cellmath__24_0_I1441 (.CO(N5034), .S(N4575), .A(N3343), .B(N4522), .CI(N4241));
ADDFX1 inst_cellmath__24_0_I1442 (.CO(N3860), .S(N3413), .A(N3957), .B(N5131), .CI(N4847));
ADDFX1 inst_cellmath__24_0_I1443 (.CO(N4764), .S(N4314), .A(N4569), .B(N3680), .CI(N3535));
ADDFXL inst_cellmath__24_0_I1444 (.CO(N3600), .S(N3144), .A(N5106), .B(N4435), .CI(N3265));
ADDFX1 inst_cellmath__24_0_I1445 (.CO(N4502), .S(N4055), .A(N5075), .B(N4168), .CI(N3904));
ADDFX1 inst_cellmath__24_0_I1446 (.CO(N3333), .S(N4953), .A(N3679), .B(N4842), .CI(N3937));
ADDFX1 inst_cellmath__24_0_I1447 (.CO(N4237), .S(N3788), .A(N3413), .B(N4575), .CI(N4804));
ADDFXL inst_cellmath__24_0_I1448 (.CO(N5138), .S(N4689), .A(N3644), .B(N4314), .CI(N4548));
ADDFX1 inst_cellmath__24_0_I1449 (.CO(N3977), .S(N3527), .A(N4055), .B(N3374), .CI(N3144));
ADDFXL inst_cellmath__24_0_I1450 (.CO(N4877), .S(N4425), .A(N4953), .B(N4281), .CI(N3788));
ADDFXL inst_cellmath__24_0_I1451 (.CO(N3710), .S(N3257), .A(N4689), .B(N3115), .CI(N4018));
ADDFXL inst_cellmath__24_0_I1452 (.CO(N4612), .S(N4159), .A(N4425), .B(N3527), .CI(N4921));
ADDFHX1 inst_cellmath__24_0_I1453 (.CO(N3447), .S(N5064), .A(N3756), .B(N3257), .CI(N4159));
ADDHX1 inst_cellmath__24_0_I1454 (.CO(N4344), .S(N3896), .A(N3874), .B(N4766));
ADDFXL inst_cellmath__24_0_I1455 (.CO(N3182), .S(N4796), .A(N4488), .B(N3303), .CI(N3592));
ADDFX1 inst_cellmath__24_0_I1456 (.CO(N4085), .S(N3633), .A(N5094), .B(N4199), .CI(N3920));
ADDFX1 inst_cellmath__24_0_I1457 (.CO(N4988), .S(N4539), .A(N4811), .B(N3639), .CI(N4534));
ADDFX1 inst_cellmath__24_0_I1458 (.CO(N3823), .S(N3365), .A(N4248), .B(N5141), .CI(N3352));
ADDFXL inst_cellmath__24_0_I1459 (.CO(N4721), .S(N4266), .A(N4858), .B(N3687), .CI(N3967));
ADDFX1 inst_cellmath__24_0_I1460 (.CO(N3553), .S(N3107), .A(N3399), .B(N4576), .CI(N4295));
ADDFHXL inst_cellmath__24_0_I1461 (.CO(N4462), .S(N4011), .A(N3494), .B(N3896), .CI(N4394));
ADDFXL inst_cellmath__24_0_I1462 (.CO(N3286), .S(N4908), .A(N3224), .B(N4129), .CI(N5034));
ADDFX1 inst_cellmath__24_0_I1463 (.CO(N4194), .S(N3747), .A(N3860), .B(N4796), .CI(N4764));
ADDFX1 inst_cellmath__24_0_I1464 (.CO(N5098), .S(N4644), .A(N4539), .B(N3633), .CI(N3365));
ADDFXL inst_cellmath__24_0_I1465 (.CO(N3929), .S(N3484), .A(N3107), .B(N4266), .CI(N3600));
ADDFX1 inst_cellmath__24_0_I1466 (.CO(N4833), .S(N4383), .A(N4502), .B(N4011), .CI(N3333));
ADDFX1 inst_cellmath__24_0_I1467 (.CO(N3671), .S(N3214), .A(N4237), .B(N4908), .CI(N3747));
ADDFXL inst_cellmath__24_0_I1468 (.CO(N4568), .S(N4120), .A(N5138), .B(N4644), .CI(N3484));
ADDFX1 inst_cellmath__24_0_I1469 (.CO(N3403), .S(N5024), .A(N4383), .B(N3977), .CI(N4877));
ADDFXL inst_cellmath__24_0_I1470 (.CO(N4304), .S(N3853), .A(N3214), .B(N4120), .CI(N3710));
ADDFHXL inst_cellmath__24_0_I1471 (.CO(N3136), .S(N4755), .A(N5024), .B(N4612), .CI(N3853));
ADDHXL inst_cellmath__24_0_I1472 (.CO(N4046), .S(N3590), .A(N3601), .B(N4775));
ADDFHXL inst_cellmath__24_0_I1473 (.CO(N4944), .S(N4494), .A(N3314), .B(N4498), .CI(N4208));
ADDFXL inst_cellmath__24_0_I1474 (.CO(N3779), .S(N3321), .A(N3930), .B(N5104), .CI(N4822));
ADDFXL inst_cellmath__24_0_I1475 (.CO(N4679), .S(N4225), .A(N4545), .B(N3649), .CI(N3362));
ADDFX1 inst_cellmath__24_0_I1476 (.CO(N3518), .S(N5127), .A(N3082), .B(N3979), .CI(N4255));
ADDFXL inst_cellmath__24_0_I1477 (.CO(N4416), .S(N3966), .A(N3694), .B(N4871), .CI(N4586));
ADDFX1 inst_cellmath__24_0_I1478 (.CO(N3248), .S(N4866), .A(N4305), .B(N3409), .CI(N3129));
ADDFXL inst_cellmath__24_0_I1479 (.CO(N4149), .S(N3699), .A(N4344), .B(N4025), .CI(N3590));
ADDFXL inst_cellmath__24_0_I1480 (.CO(N5054), .S(N4603), .A(N4085), .B(N3182), .CI(N4988));
ADDFXL inst_cellmath__24_0_I1481 (.CO(N3888), .S(N3437), .A(N4721), .B(N3823), .CI(N3553));
ADDFXL inst_cellmath__24_0_I1482 (.CO(N4786), .S(N4334), .A(N4494), .B(N3321), .CI(N4225));
ADDFX1 inst_cellmath__24_0_I1483 (.CO(N3625), .S(N3171), .A(N5127), .B(N3966), .CI(N4866));
ADDFXL inst_cellmath__24_0_I1484 (.CO(N4529), .S(N4074), .A(N3286), .B(N4462), .CI(N3699));
ADDFHX1 inst_cellmath__24_0_I1485 (.CO(N3355), .S(N4979), .A(N3437), .B(N4194), .CI(N4603));
ADDFX1 inst_cellmath__24_0_I1486 (.CO(N4257), .S(N3813), .A(N3929), .B(N5098), .CI(N4334));
ADDFXL inst_cellmath__24_0_I1487 (.CO(N3096), .S(N4710), .A(N4833), .B(N3171), .CI(N4074));
ADDFXL inst_cellmath__24_0_I1488 (.CO(N4000), .S(N3546), .A(N4979), .B(N3671), .CI(N4568));
ADDFXL inst_cellmath__24_0_I1489 (.CO(N4900), .S(N4452), .A(N4710), .B(N3813), .CI(N3403));
ADDFXL inst_cellmath__24_0_I1490 (.CO(N3736), .S(N3278), .A(N3546), .B(N4304), .CI(N4452));
ADDHX1 inst_cellmath__24_0_I1491 (.CO(N4634), .S(N4180), .A(N3612), .B(N4506));
ADDFHXL inst_cellmath__24_0_I1492 (.CO(N3472), .S(N5088), .A(N4217), .B(N3323), .CI(N5111));
ADDFXL inst_cellmath__24_0_I1493 (.CO(N4373), .S(N3922), .A(N3659), .B(N3938), .CI(N4829));
ADDFX1 inst_cellmath__24_0_I1494 (.CO(N3205), .S(N4821), .A(N4553), .B(N3372), .CI(N4263));
ADDFHX1 inst_cellmath__24_0_I1495 (.CO(N4109), .S(N3661), .A(N3988), .B(N3091), .CI(N4880));
ADDFXL inst_cellmath__24_0_I1496 (.CO(N5014), .S(N4563), .A(N4595), .B(N3703), .CI(N3419));
ADDFX1 inst_cellmath__24_0_I1497 (.CO(N3846), .S(N3393), .A(N3137), .B(N4315), .CI(N4035));
ADDFXL inst_cellmath__24_0_I1498 (.CO(N4744), .S(N4298), .A(N4926), .B(N3754), .CI(N4046));
ADDFX1 inst_cellmath__24_0_I1499 (.CO(N3581), .S(N3128), .A(N4180), .B(N4944), .CI(N3779));
ADDFXL inst_cellmath__24_0_I1500 (.CO(N4487), .S(N4034), .A(N4679), .B(N3518), .CI(N4416));
ADDFXL inst_cellmath__24_0_I1501 (.CO(N3311), .S(N4937), .A(N3248), .B(N5088), .CI(N3922));
ADDFXL inst_cellmath__24_0_I1502 (.CO(N4215), .S(N3772), .A(N4821), .B(N3661), .CI(N4563));
ADDFX1 inst_cellmath__24_0_I1503 (.CO(N5119), .S(N4670), .A(N4149), .B(N3393), .CI(N5054));
ADDFHXL inst_cellmath__24_0_I1504 (.CO(N3955), .S(N3510), .A(N3888), .B(N4298), .CI(N4786));
ADDFX1 inst_cellmath__24_0_I1505 (.CO(N4856), .S(N4408), .A(N4034), .B(N3625), .CI(N3128));
ADDFHXL inst_cellmath__24_0_I1506 (.CO(N3691), .S(N3239), .A(N3772), .B(N4937), .CI(N4529));
ADDFHXL inst_cellmath__24_0_I1507 (.CO(N4592), .S(N4140), .A(N3355), .B(N4670), .CI(N3510));
ADDFHXL inst_cellmath__24_0_I1508 (.CO(N3426), .S(N5046), .A(N4408), .B(N4257), .CI(N3239));
ADDFXL inst_cellmath__24_0_I1509 (.CO(N4327), .S(N3877), .A(N4140), .B(N3096), .CI(N4000));
ADDHX1 inst_cellmath__24_0_I1511 (.CO(N4065), .S(N3616), .A(N4515), .B(N3335));
ADDFHXL inst_cellmath__24_0_I1512 (.CO(N4969), .S(N4519), .A(N3947), .B(N4228), .CI(N5120));
ADDFHX1 inst_cellmath__24_0_I1513 (.CO(N3804), .S(N3347), .A(N4839), .B(N3668), .CI(N4561));
ADDFHXL inst_cellmath__24_0_I1514 (.CO(N4702), .S(N4249), .A(N4275), .B(N3100), .CI(N3384));
ADDFXL inst_cellmath__24_0_I1515 (.CO(N3538), .S(N3086), .A(N4890), .B(N3996), .CI(N3714));
ADDFXL inst_cellmath__24_0_I1516 (.CO(N4444), .S(N3991), .A(N3430), .B(N4323), .CI(N4604));
ADDFXL inst_cellmath__24_0_I1517 (.CO(N3270), .S(N4892), .A(N4042), .B(N4938), .CI(N3145));
ADDFX1 inst_cellmath__24_0_I1518 (.CO(N4172), .S(N3728), .A(N4649), .B(N3762), .CI(N3477));
ADDFHXL inst_cellmath__24_0_I1519 (.CO(N5080), .S(N4625), .A(N3616), .B(N4634), .CI(N3472));
ADDFHXL inst_cellmath__24_0_I1520 (.CO(N3912), .S(N3463), .A(N4109), .B(N3205), .CI(N4373));
ADDFHXL inst_cellmath__24_0_I1521 (.CO(N4810), .S(N4363), .A(N3846), .B(N5014), .CI(N4519));
ADDFXL inst_cellmath__24_0_I1522 (.CO(N3650), .S(N3195), .A(N3347), .B(N4249), .CI(N4744));
ADDFX1 inst_cellmath__24_0_I1523 (.CO(N4554), .S(N4099), .A(N3991), .B(N3086), .CI(N4892));
ADDFX1 inst_cellmath__24_0_I1524 (.CO(N3383), .S(N5004), .A(N3581), .B(N3728), .CI(N4487));
ADDFXL inst_cellmath__24_0_I1525 (.CO(N4287), .S(N3836), .A(N3463), .B(N4625), .CI(N3311));
ADDFX1 inst_cellmath__24_0_I1526 (.CO(N3121), .S(N4733), .A(N4363), .B(N4215), .CI(N3195));
ADDFX1 inst_cellmath__24_0_I1527 (.CO(N4024), .S(N3571), .A(N4099), .B(N5119), .CI(N3955));
ADDFXL inst_cellmath__24_0_I1528 (.CO(N4928), .S(N4478), .A(N5004), .B(N4856), .CI(N3836));
ADDFHXL inst_cellmath__24_0_I1529 (.CO(N3761), .S(N3300), .A(N4733), .B(N3691), .CI(N4592));
ADDFHXL inst_cellmath__24_0_I1530 (.CO(N4658), .S(N4207), .A(N4478), .B(N3571), .CI(N3426));
ADDHX1 inst_cellmath__24_0_I1532 (.CO(N4401), .S(N3944), .A(N3468), .B(N4238));
ADDFXL inst_cellmath__24_0_I1533 (.CO(N3229), .S(N4846), .A(N3344), .B(N5132), .CI(N3958));
ADDFHX1 inst_cellmath__24_0_I1534 (.CO(N4134), .S(N3683), .A(N4570), .B(N3677), .CI(N4848));
ADDFHX1 inst_cellmath__24_0_I1535 (.CO(N5038), .S(N4582), .A(N3112), .B(N3394), .CI(N4285));
ADDFXL inst_cellmath__24_0_I1536 (.CO(N3868), .S(N3417), .A(N4898), .B(N4008), .CI(N3724));
ADDFXL inst_cellmath__24_0_I1537 (.CO(N4769), .S(N4319), .A(N3441), .B(N4613), .CI(N4330));
ADDFX1 inst_cellmath__24_0_I1538 (.CO(N3607), .S(N3152), .A(N4051), .B(N3154), .CI(N4945));
ADDFX1 inst_cellmath__24_0_I1539 (.CO(N4510), .S(N4058), .A(N4659), .B(N3773), .CI(N3489));
ADDFXL inst_cellmath__24_0_I1540 (.CO(N3339), .S(N4959), .A(N4065), .B(N4380), .CI(N3944));
ADDFHXL inst_cellmath__24_0_I1541 (.CO(N4242), .S(N3795), .A(N3804), .B(N4702), .CI(N4969));
ADDFXL inst_cellmath__24_0_I1542 (.CO(N5145), .S(N4693), .A(N4444), .B(N3270), .CI(N3538));
ADDFX1 inst_cellmath__24_0_I1543 (.CO(N3982), .S(N3532), .A(N4846), .B(N4172), .CI(N3683));
ADDFX1 inst_cellmath__24_0_I1544 (.CO(N4882), .S(N4433), .A(N3417), .B(N4582), .CI(N4319));
ADDFHXL inst_cellmath__24_0_I1545 (.CO(N3717), .S(N3262), .A(N4058), .B(N3152), .CI(N3912));
ADDFHX1 inst_cellmath__24_0_I1546 (.CO(N4617), .S(N4164), .A(N5080), .B(N4810), .CI(N4959));
ADDFXL inst_cellmath__24_0_I1547 (.CO(N3452), .S(N5070), .A(N3650), .B(N3795), .CI(N4693));
ADDFXL inst_cellmath__24_0_I1548 (.CO(N4352), .S(N3901), .A(N3532), .B(N4554), .CI(N4433));
ADDFXL inst_cellmath__24_0_I1549 (.CO(N3186), .S(N4802), .A(N3383), .B(N3262), .CI(N4287));
ADDFHXL inst_cellmath__24_0_I1550 (.CO(N4089), .S(N3640), .A(N3121), .B(N4164), .CI(N5070));
ADDFXL inst_cellmath__24_0_I1551 (.CO(N4995), .S(N4546), .A(N3901), .B(N4024), .CI(N4802));
ADDFHXL inst_cellmath__24_0_I1552 (.CO(N3828), .S(N3370), .A(N3640), .B(N4928), .CI(N3761));
ADDHX1 inst_cellmath__24_0_I1554 (.CO(N3562), .S(N3113), .A(N4371), .B(N3968));
ADDFXL inst_cellmath__24_0_I1555 (.CO(N4467), .S(N4016), .A(N5142), .B(N3684), .CI(N4859));
ADDFXL inst_cellmath__24_0_I1556 (.CO(N3291), .S(N4917), .A(N4577), .B(N3400), .CI(N4296));
ADDFXL inst_cellmath__24_0_I1557 (.CO(N4198), .S(N3753), .A(N4017), .B(N3120), .CI(N4905));
ADDFHXL inst_cellmath__24_0_I1558 (.CO(N5102), .S(N4648), .A(N4622), .B(N3732), .CI(N3451));
ADDFXL inst_cellmath__24_0_I1559 (.CO(N3936), .S(N3491), .A(N4059), .B(N3162), .CI(N4338));
ADDFXL inst_cellmath__24_0_I1560 (.CO(N4836), .S(N4390), .A(N4954), .B(N3780), .CI(N4667));
ADDFX1 inst_cellmath__24_0_I1561 (.CO(N3675), .S(N3221), .A(N4391), .B(N3500), .CI(N3211));
ADDFHXL inst_cellmath__24_0_I1562 (.CO(N4574), .S(N4126), .A(N3113), .B(N4401), .CI(N3229));
ADDFHXL inst_cellmath__24_0_I1563 (.CO(N3407), .S(N5030), .A(N5038), .B(N4134), .CI(N3868));
ADDFHXL inst_cellmath__24_0_I1564 (.CO(N4311), .S(N3858), .A(N3607), .B(N4510), .CI(N4769));
ADDFXL inst_cellmath__24_0_I1565 (.CO(N3142), .S(N4761), .A(N3753), .B(N4016), .CI(N4917));
ADDFX1 inst_cellmath__24_0_I1566 (.CO(N4049), .S(N3596), .A(N4648), .B(N4390), .CI(N3491));
ADDFXL inst_cellmath__24_0_I1567 (.CO(N4950), .S(N4500), .A(N3339), .B(N3221), .CI(N4242));
ADDFHXL inst_cellmath__24_0_I1568 (.CO(N3785), .S(N3327), .A(N5145), .B(N4126), .CI(N5030));
ADDFHXL inst_cellmath__24_0_I1569 (.CO(N4684), .S(N4233), .A(N3858), .B(N3982), .CI(N4882));
ADDFX1 inst_cellmath__24_0_I1570 (.CO(N3524), .S(N5134), .A(N4761), .B(N3717), .CI(N3596));
ADDFHXL inst_cellmath__24_0_I1571 (.CO(N4421), .S(N3972), .A(N4617), .B(N4500), .CI(N3452));
ADDFHX1 inst_cellmath__24_0_I1572 (.CO(N3253), .S(N4872), .A(N4233), .B(N3327), .CI(N4352));
ADDFHXL inst_cellmath__24_0_I1573 (.CO(N4155), .S(N3706), .A(N5134), .B(N3186), .CI(N3972));
ADDFHXL inst_cellmath__24_0_I1574 (.CO(N5060), .S(N4608), .A(N4872), .B(N4089), .CI(N4995));
ADDFHXL inst_cellmath__24_0_I1575 (.CO(N3892), .S(N3442), .A(N3828), .B(N3706), .CI(N4608));
ADDFXL inst_cellmath__24_0_I1576 (.CO(N4792), .S(N4342), .A(N4868), .B(N3201), .CI(N3695));
ADDFHXL inst_cellmath__24_0_I1577 (.CO(N3631), .S(N3177), .A(N3410), .B(N4587), .CI(N4302));
ADDFXL inst_cellmath__24_0_I1578 (.CO(N4535), .S(N4080), .A(N4026), .B(N4916), .CI(N3130));
ADDFX1 inst_cellmath__24_0_I1579 (.CO(N3361), .S(N4986), .A(N4633), .B(N3742), .CI(N3461));
ADDFX1 inst_cellmath__24_0_I1580 (.CO(N4265), .S(N3817), .A(N4348), .B(N3172), .CI(N4069));
ADDFX1 inst_cellmath__24_0_I1581 (.CO(N3101), .S(N4716), .A(N3789), .B(N4964), .CI(N4676));
ADDFX1 inst_cellmath__24_0_I1582 (.CO(N4007), .S(N3552), .A(N4402), .B(N11813), .CI(N3222));
ADDFXL inst_cellmath__24_0_I1583 (.CO(N4907), .S(N4457), .A(N3562), .B(N4113), .CI(N4467));
ADDFXL inst_cellmath__24_0_I1584 (.CO(N3743), .S(N3283), .A(N4198), .B(N5102), .CI(N3291));
ADDFXL inst_cellmath__24_0_I1585 (.CO(N4639), .S(N4188), .A(N4836), .B(N3936), .CI(N3675));
ADDFHXL inst_cellmath__24_0_I1586 (.CO(N3480), .S(N5092), .A(N4342), .B(N4080), .CI(N3177));
ADDFXL inst_cellmath__24_0_I1587 (.CO(N4379), .S(N3927), .A(N3817), .B(N4716), .CI(N4986));
ADDFHXL inst_cellmath__24_0_I1588 (.CO(N3210), .S(N4828), .A(N4574), .B(N3552), .CI(N3407));
ADDFX1 inst_cellmath__24_0_I1589 (.CO(N4115), .S(N3667), .A(N4311), .B(N4457), .CI(N3142));
ADDFXL inst_cellmath__24_0_I1590 (.CO(N5020), .S(N4566), .A(N4049), .B(N3283), .CI(N4188));
ADDFX1 inst_cellmath__24_0_I1591 (.CO(N3850), .S(N3398), .A(N4950), .B(N5092), .CI(N3927));
ADDFHXL inst_cellmath__24_0_I1592 (.CO(N4752), .S(N4301), .A(N4828), .B(N3785), .CI(N4684));
ADDFXL inst_cellmath__24_0_I1593 (.CO(N3586), .S(N3134), .A(N4566), .B(N3667), .CI(N3524));
ADDFHXL inst_cellmath__24_0_I1594 (.CO(N4492), .S(N4041), .A(N3398), .B(N4421), .CI(N4301));
ADDFHXL inst_cellmath__24_0_I1595 (.CO(N3318), .S(N4941), .A(N3134), .B(N3253), .CI(N4155));
ADDFHXL inst_cellmath__24_0_I1596 (.CO(N4221), .S(N3777), .A(N5060), .B(N4041), .CI(N4941));
ADDFHXL inst_cellmath__24_0_I1597 (.CO(N5124), .S(N4675), .A(N4104), .B(N4596), .CI(N3420));
ADDFXL inst_cellmath__24_0_I1598 (.CO(N3963), .S(N3515), .A(N3138), .B(N4312), .CI(N4036));
ADDFXL inst_cellmath__24_0_I1599 (.CO(N4863), .S(N4413), .A(N4927), .B(N3752), .CI(N4640));
ADDFX1 inst_cellmath__24_0_I1600 (.CO(N3696), .S(N3244), .A(N4359), .B(N3183), .CI(N3469));
ADDFXL inst_cellmath__24_0_I1601 (.CO(N4600), .S(N4147), .A(N4079), .B(N4973), .CI(N3797));
ADDFX1 inst_cellmath__24_0_I1602 (.CO(N3432), .S(N5051), .A(N4685), .B(N3519), .CI(N4409));
ADDFX1 inst_cellmath__24_0_I1603 (.CO(N4331), .S(N3884), .A(N4124), .B(N3230), .CI(N5021));
ADDFHXL inst_cellmath__24_0_I1604 (.CO(N3167), .S(N4784), .A(N4535), .B(N4792), .CI(N3631));
ADDFHXL inst_cellmath__24_0_I1605 (.CO(N4071), .S(N3622), .A(N4265), .B(N3361), .CI(N3101));
ADDFX1 inst_cellmath__24_0_I1606 (.CO(N4976), .S(N4525), .A(N3515), .B(N4007), .CI(N4675));
ADDFXL inst_cellmath__24_0_I1607 (.CO(N3810), .S(N3354), .A(N4413), .B(N3244), .CI(N4147));
ADDFXL inst_cellmath__24_0_I1608 (.CO(N4707), .S(N4254), .A(N3884), .B(N5051), .CI(N4907));
ADDFHXL inst_cellmath__24_0_I1609 (.CO(N3543), .S(N3093), .A(N4639), .B(N3743), .CI(N3480));
ADDFX1 inst_cellmath__24_0_I1610 (.CO(N4450), .S(N3998), .A(N4784), .B(N3622), .CI(N4379));
ADDFX1 inst_cellmath__24_0_I1611 (.CO(N3276), .S(N4897), .A(N3210), .B(N4525), .CI(N3354));
ADDFHXL inst_cellmath__24_0_I1612 (.CO(N4177), .S(N3734), .A(N4115), .B(N4254), .CI(N5020));
ADDFHXL inst_cellmath__24_0_I1613 (.CO(N5086), .S(N4632), .A(N3093), .B(N3850), .CI(N3998));
ADDFHXL inst_cellmath__24_0_I1614 (.CO(N3918), .S(N3471), .A(N4897), .B(N4752), .CI(N3734));
ADDFHXL inst_cellmath__24_0_I1615 (.CO(N4819), .S(N4370), .A(N4632), .B(N3586), .CI(N4492));
ADDFHXL inst_cellmath__24_0_I1616 (.CO(N3658), .S(N3200), .A(N3318), .B(N3471), .CI(N4370));
ADDFXL inst_cellmath__24_0_I1617 (.CO(N4559), .S(N4107), .A(N5012), .B(N3146), .CI(N4320));
ADDFXL inst_cellmath__24_0_I1618 (.CO(N3392), .S(N5011), .A(N4043), .B(N4935), .CI(N3760));
ADDFXL inst_cellmath__24_0_I1619 (.CO(N4294), .S(N3841), .A(N4368), .B(N3478), .CI(N4650));
ADDFXL inst_cellmath__24_0_I1620 (.CO(N3125), .S(N4743), .A(N4982), .B(N3191), .CI(N4088));
ADDFXL inst_cellmath__24_0_I1621 (.CO(N4033), .S(N3578), .A(N3528), .B(N4695), .CI(N3805));
ADDFXL inst_cellmath__24_0_I1622 (.CO(N4934), .S(N4482), .A(N3238), .B(N4417), .CI(N4133));
ADDFHXL inst_cellmath__24_0_I1623 (.CO(N3768), .S(N3309), .A(N3851), .B(N5031), .CI(N5124));
ADDFXL inst_cellmath__24_0_I1624 (.CO(N4666), .S(N4212), .A(N4863), .B(N3963), .CI(N3696));
ADDFX1 inst_cellmath__24_0_I1625 (.CO(N3507), .S(N5115), .A(N3432), .B(N4600), .CI(N4331));
ADDFXL inst_cellmath__24_0_I1626 (.CO(N4406), .S(N3953), .A(N4107), .B(N5011), .CI(N3841));
ADDFXL inst_cellmath__24_0_I1627 (.CO(N3237), .S(N4853), .A(N3578), .B(N4743), .CI(N4482));
ADDFHXL inst_cellmath__24_0_I1628 (.CO(N4139), .S(N3688), .A(N4071), .B(N3167), .CI(N3309));
ADDFXL inst_cellmath__24_0_I1629 (.CO(N5043), .S(N4591), .A(N4212), .B(N4976), .CI(N3810));
ADDFXL inst_cellmath__24_0_I1630 (.CO(N3875), .S(N3424), .A(N4707), .B(N5115), .CI(N3953));
ADDFHXL inst_cellmath__24_0_I1631 (.CO(N4777), .S(N4325), .A(N4853), .B(N3543), .CI(N4450));
ADDFXL inst_cellmath__24_0_I1632 (.CO(N3613), .S(N3159), .A(N4591), .B(N3688), .CI(N3276));
ADDFHXL inst_cellmath__24_0_I1633 (.CO(N4517), .S(N4062), .A(N3424), .B(N4177), .CI(N4325));
ADDFHXL inst_cellmath__24_0_I1634 (.CO(N3345), .S(N4966), .A(N3159), .B(N5086), .CI(N3918));
ADDFHXL inst_cellmath__24_0_I1635 (.CO(N4247), .S(N3802), .A(N4819), .B(N4062), .CI(N4966));
ADDFX1 inst_cellmath__24_0_I1636 (.CO(N3084), .S(N4699), .A(N4052), .B(N3842), .CI(N4942));
ADDFXL inst_cellmath__24_0_I1637 (.CO(N3990), .S(N3537), .A(N4660), .B(N3774), .CI(N3490));
ADDFXL inst_cellmath__24_0_I1638 (.CO(N4888), .S(N4442), .A(N4098), .B(N3202), .CI(N4378));
ADDFXL inst_cellmath__24_0_I1639 (.CO(N3726), .S(N3267), .A(N3814), .B(N4993), .CI(N4705));
ADDFXL inst_cellmath__24_0_I1640 (.CO(N4623), .S(N4170), .A(N3245), .B(N3536), .CI(N4426));
ADDFX1 inst_cellmath__24_0_I1641 (.CO(N3459), .S(N5078), .A(N5039), .B(N4141), .CI(N3859));
ADDFX1 inst_cellmath__24_0_I1642 (.CO(N4361), .S(N3909), .A(N4750), .B(N3392), .CI(N4559));
ADDFX1 inst_cellmath__24_0_I1643 (.CO(N3193), .S(N4808), .A(N3125), .B(N4033), .CI(N4294));
ADDFXL inst_cellmath__24_0_I1644 (.CO(N4096), .S(N3647), .A(N4934), .B(N4699), .CI(N3537));
ADDFXL inst_cellmath__24_0_I1645 (.CO(N5003), .S(N4551), .A(N4170), .B(N4442), .CI(N3267));
ADDFHXL inst_cellmath__24_0_I1646 (.CO(N3833), .S(N3379), .A(N5078), .B(N3768), .CI(N4666));
ADDFXL inst_cellmath__24_0_I1647 (.CO(N4729), .S(N4284), .A(N3909), .B(N3507), .CI(N4808));
ADDFX1 inst_cellmath__24_0_I1648 (.CO(N3570), .S(N3118), .A(N3237), .B(N4406), .CI(N3647));
ADDFHXL inst_cellmath__24_0_I1649 (.CO(N4474), .S(N4020), .A(N4551), .B(N4139), .CI(N3379));
ADDFXL inst_cellmath__24_0_I1650 (.CO(N3296), .S(N4924), .A(N5043), .B(N3875), .CI(N4284));
ADDFHXL inst_cellmath__24_0_I1651 (.CO(N4205), .S(N3758), .A(N4777), .B(N3118), .CI(N4020));
ADDFHXL inst_cellmath__24_0_I1652 (.CO(N5107), .S(N4657), .A(N4924), .B(N3613), .CI(N4517));
ADDFHXL inst_cellmath__24_0_I1653 (.CO(N3943), .S(N3498), .A(N3345), .B(N3758), .CI(N4657));
ADDFX1 inst_cellmath__24_0_I1654 (.CO(N4843), .S(N4397), .A(N3781), .B(N4740), .CI(N4668));
ADDFXL inst_cellmath__24_0_I1655 (.CO(N3681), .S(N3228), .A(N4389), .B(N3501), .CI(N3212));
ADDFXL inst_cellmath__24_0_I1656 (.CO(N4581), .S(N4131), .A(N5001), .B(N4105), .CI(N3824));
ADDFXL inst_cellmath__24_0_I1657 (.CO(N3415), .S(N5036), .A(N4714), .B(N3541), .CI(N4436));
ADDFXL inst_cellmath__24_0_I1658 (.CO(N4316), .S(N3867), .A(N4150), .B(N3254), .CI(N5047));
ADDFXL inst_cellmath__24_0_I1659 (.CO(N3150), .S(N4767), .A(N4760), .B(N3869), .CI(N3587));
ADDFX1 inst_cellmath__24_0_I1660 (.CO(N4056), .S(N3602), .A(N3084), .B(N4888), .CI(N3990));
ADDFX1 inst_cellmath__24_0_I1661 (.CO(N4956), .S(N4507), .A(N4623), .B(N3726), .CI(N3459));
ADDFX1 inst_cellmath__24_0_I1662 (.CO(N3793), .S(N3337), .A(N3228), .B(N4397), .CI(N4131));
ADDFXL inst_cellmath__24_0_I1663 (.CO(N4690), .S(N4239), .A(N3867), .B(N4767), .CI(N5036));
ADDFX1 inst_cellmath__24_0_I1664 (.CO(N3529), .S(N5143), .A(N3193), .B(N4361), .CI(N4096));
ADDFX1 inst_cellmath__24_0_I1665 (.CO(N4431), .S(N3980), .A(N3602), .B(N5003), .CI(N4507));
ADDFXL inst_cellmath__24_0_I1666 (.CO(N3258), .S(N4878), .A(N3833), .B(N4239), .CI(N3337));
ADDFXL inst_cellmath__24_0_I1667 (.CO(N4161), .S(N3715), .A(N4729), .B(N3570), .CI(N5143));
ADDFX1 inst_cellmath__24_0_I1668 (.CO(N5068), .S(N4615), .A(N4474), .B(N3980), .CI(N4878));
ADDFHXL inst_cellmath__24_0_I1669 (.CO(N3898), .S(N3449), .A(N3715), .B(N3296), .CI(N4205));
ADDFHXL inst_cellmath__24_0_I1670 (.CO(N4799), .S(N4350), .A(N5107), .B(N4615), .CI(N3449));
ADDFXL inst_cellmath__24_0_I1671 (.CO(N3638), .S(N3184), .A(N3508), .B(N3579), .CI(N4400));
ADDFXL inst_cellmath__24_0_I1672 (.CO(N4543), .S(N4086), .A(N5009), .B(N4114), .CI(N3223));
ADDFXL inst_cellmath__24_0_I1673 (.CO(N3368), .S(N4994), .A(N4724), .B(N3832), .CI(N3549));
ADDFX1 inst_cellmath__24_0_I1674 (.CO(N4274), .S(N3825), .A(N3263), .B(N4160), .CI(N4445));
ADDFX1 inst_cellmath__24_0_I1675 (.CO(N3110), .S(N4722), .A(N3876), .B(N5055), .CI(N4770));
ADDFX1 inst_cellmath__24_0_I1676 (.CO(N4014), .S(N3561), .A(N4493), .B(N3597), .CI(N4843));
ADDFX1 inst_cellmath__24_0_I1677 (.CO(N4915), .S(N4465), .A(N4581), .B(N3681), .CI(N3415));
ADDFX1 inst_cellmath__24_0_I1678 (.CO(N3749), .S(N3288), .A(N3150), .B(N4316), .CI(N3184));
ADDFX1 inst_cellmath__24_0_I1679 (.CO(N4646), .S(N4197), .A(N4994), .B(N4086), .CI(N3825));
ADDFX1 inst_cellmath__24_0_I1680 (.CO(N3488), .S(N5100), .A(N4056), .B(N4722), .CI(N4956));
ADDFX1 inst_cellmath__24_0_I1681 (.CO(N4386), .S(N3933), .A(N3793), .B(N3561), .CI(N4465));
ADDFHXL inst_cellmath__24_0_I1682 (.CO(N3217), .S(N4835), .A(N3288), .B(N4690), .CI(N4197));
ADDFX1 inst_cellmath__24_0_I1683 (.CO(N4123), .S(N3673), .A(N4431), .B(N3529), .CI(N5100));
ADDFX1 inst_cellmath__24_0_I1684 (.CO(N5027), .S(N4572), .A(N3933), .B(N3258), .CI(N4835));
ADDFHXL inst_cellmath__24_0_I1685 (.CO(N3855), .S(N3406), .A(N3673), .B(N4161), .CI(N5068));
ADDFHXL inst_cellmath__24_0_I1686 (.CO(N4759), .S(N4307), .A(N3898), .B(N4572), .CI(N3406));
ADDFX1 inst_cellmath__24_0_I1687 (.CO(N3593), .S(N3140), .A(N3231), .B(N4483), .CI(N4125));
ADDFXL inst_cellmath__24_0_I1688 (.CO(N4499), .S(N4047), .A(N3843), .B(N5019), .CI(N4731));
ADDFXL inst_cellmath__24_0_I1689 (.CO(N3324), .S(N4948), .A(N4453), .B(N3559), .CI(N3273));
ADDFX1 inst_cellmath__24_0_I1690 (.CO(N4229), .S(N3784), .A(N5065), .B(N4169), .CI(N3885));
ADDFX1 inst_cellmath__24_0_I1691 (.CO(N5133), .S(N4681), .A(N3608), .B(N4779), .CI(N4501));
ADDFX1 inst_cellmath__24_0_I1692 (.CO(N3969), .S(N3521), .A(N3638), .B(N3317), .CI(N4543));
ADDFX1 inst_cellmath__24_0_I1693 (.CO(N4869), .S(N4420), .A(N4274), .B(N3368), .CI(N3110));
ADDFXL inst_cellmath__24_0_I1694 (.CO(N3705), .S(N3250), .A(N4948), .B(N3140), .CI(N4047));
ADDFX1 inst_cellmath__24_0_I1695 (.CO(N4605), .S(N4153), .A(N4681), .B(N3784), .CI(N4014));
ADDFX1 inst_cellmath__24_0_I1696 (.CO(N3439), .S(N5059), .A(N3749), .B(N4915), .CI(N3521));
ADDFXL inst_cellmath__24_0_I1697 (.CO(N4339), .S(N3889), .A(N4420), .B(N4646), .CI(N3250));
ADDFX1 inst_cellmath__24_0_I1698 (.CO(N3174), .S(N4789), .A(N4153), .B(N3488), .CI(N4386));
ADDFX1 inst_cellmath__24_0_I1699 (.CO(N4077), .S(N3628), .A(N3217), .B(N5059), .CI(N3889));
ADDFHXL inst_cellmath__24_0_I1700 (.CO(N4983), .S(N4532), .A(N4123), .B(N4789), .CI(N5027));
ADDFHXL inst_cellmath__24_0_I1701 (.CO(N3815), .S(N3359), .A(N3628), .B(N3855), .CI(N4532));
ADDFX1 inst_cellmath__24_0_I1702 (.CO(N4712), .S(N4262), .A(N5029), .B(N3307), .CI(N3852));
ADDFX1 inst_cellmath__24_0_I1703 (.CO(N3550), .S(N3098), .A(N4741), .B(N3569), .CI(N4464));
ADDFX1 inst_cellmath__24_0_I1704 (.CO(N4455), .S(N4004), .A(N5071), .B(N3282), .CI(N4175));
ADDFX1 inst_cellmath__24_0_I1705 (.CO(N3280), .S(N4904), .A(N4787), .B(N3893), .CI(N3617));
ADDFX1 inst_cellmath__24_0_I1706 (.CO(N4186), .S(N3740), .A(N3326), .B(N4508), .CI(N4222));
ADDFX1 inst_cellmath__24_0_I1707 (.CO(N5090), .S(N4637), .A(N4499), .B(N3593), .CI(N3324));
ADDFX1 inst_cellmath__24_0_I1708 (.CO(N3924), .S(N3476), .A(N5133), .B(N4229), .CI(N4262));
ADDFX1 inst_cellmath__24_0_I1709 (.CO(N4826), .S(N4376), .A(N4004), .B(N4904), .CI(N3098));
ADDFX1 inst_cellmath__24_0_I1710 (.CO(N3664), .S(N3207), .A(N3969), .B(N3740), .CI(N4869));
ADDFXL inst_cellmath__24_0_I1711 (.CO(N4564), .S(N4112), .A(N4637), .B(N3705), .CI(N4605));
ADDFX1 inst_cellmath__24_0_I1712 (.CO(N3397), .S(N5017), .A(N4376), .B(N3476), .CI(N3439));
ADDFX1 inst_cellmath__24_0_I1713 (.CO(N4299), .S(N3848), .A(N4339), .B(N3207), .CI(N4112));
ADDFHXL inst_cellmath__24_0_I1714 (.CO(N3131), .S(N4749), .A(N5017), .B(N3174), .CI(N4077));
ADDFHXL inst_cellmath__24_0_I1715 (.CO(N4039), .S(N3584), .A(N4983), .B(N3848), .CI(N4749));
ADDFX1 inst_cellmath__24_0_I1716 (.CO(N4939), .S(N4489), .A(N4751), .B(N4213), .CI(N3576));
ADDFXL inst_cellmath__24_0_I1717 (.CO(N3775), .S(N3316), .A(N4183), .B(N4476), .CI(N3290));
ADDFX1 inst_cellmath__24_0_I1718 (.CO(N4673), .S(N4219), .A(N3905), .B(N5081), .CI(N4797));
ADDFX1 inst_cellmath__24_0_I1719 (.CO(N3512), .S(N5121), .A(N4518), .B(N3626), .CI(N3340));
ADDFX1 inst_cellmath__24_0_I1720 (.CO(N4410), .S(N3960), .A(N5125), .B(N4234), .CI(N4712));
ADDFX1 inst_cellmath__24_0_I1721 (.CO(N3241), .S(N4860), .A(N4455), .B(N3550), .CI(N3280));
ADDFX1 inst_cellmath__24_0_I1722 (.CO(N4142), .S(N3692), .A(N4489), .B(N4186), .CI(N3316));
ADDFX1 inst_cellmath__24_0_I1723 (.CO(N5049), .S(N4597), .A(N5121), .B(N4219), .CI(N5090));
ADDFXL inst_cellmath__24_0_I1724 (.CO(N3881), .S(N3428), .A(N3960), .B(N3924), .CI(N4826));
ADDFX1 inst_cellmath__24_0_I1725 (.CO(N4780), .S(N4328), .A(N3692), .B(N4860), .CI(N3664));
ADDFX1 inst_cellmath__24_0_I1726 (.CO(N3621), .S(N3163), .A(N4564), .B(N4597), .CI(N3428));
ADDFX1 inst_cellmath__24_0_I1727 (.CO(N4520), .S(N4067), .A(N4328), .B(N3397), .CI(N4299));
ADDFHXL inst_cellmath__24_0_I1728 (.CO(N3350), .S(N4974), .A(N3131), .B(N3163), .CI(N4067));
ADDFX1 inst_cellmath__24_0_I1729 (.CO(N4253), .S(N3806), .A(N4484), .B(N5116), .CI(N3298));
ADDFX1 inst_cellmath__24_0_I1730 (.CO(N3088), .S(N4703), .A(N5089), .B(N4196), .CI(N3915));
ADDFX1 inst_cellmath__24_0_I1731 (.CO(N3994), .S(N3542), .A(N3634), .B(N4805), .CI(N4526));
ADDFX1 inst_cellmath__24_0_I1732 (.CO(N4896), .S(N4446), .A(N4243), .B(N3348), .CI(N5135));
ADDFX1 inst_cellmath__24_0_I1733 (.CO(N3730), .S(N3271), .A(N4939), .B(N3961), .CI(N3775));
ADDFX1 inst_cellmath__24_0_I1734 (.CO(N4628), .S(N4176), .A(N3512), .B(N4673), .CI(N3806));
ADDFX1 inst_cellmath__24_0_I1735 (.CO(N3467), .S(N5082), .A(N3542), .B(N4703), .CI(N4446));
ADDFXL inst_cellmath__24_0_I1736 (.CO(N4366), .S(N3913), .A(N3241), .B(N4410), .CI(N4142));
ADDFX1 inst_cellmath__24_0_I1737 (.CO(N3197), .S(N4816), .A(N4176), .B(N3271), .CI(N5049));
ADDFX1 inst_cellmath__24_0_I1738 (.CO(N4103), .S(N3653), .A(N3881), .B(N5082), .CI(N3913));
ADDFX1 inst_cellmath__24_0_I1739 (.CO(N5006), .S(N4555), .A(N4816), .B(N4780), .CI(N3621));
ADDFX1 inst_cellmath__24_0_I1740 (.CO(N3839), .S(N3388), .A(N4520), .B(N3653), .CI(N4555));
ADDFX1 inst_cellmath__24_0_I1741 (.CO(N4739), .S(N4289), .A(N4203), .B(N3951), .CI(N5099));
ADDFX1 inst_cellmath__24_0_I1742 (.CO(N3574), .S(N3122), .A(N4814), .B(N3926), .CI(N3641));
ADDFX1 inst_cellmath__24_0_I1743 (.CO(N4480), .S(N4030), .A(N3356), .B(N4536), .CI(N4250));
ADDFX1 inst_cellmath__24_0_I1744 (.CO(N3306), .S(N4929), .A(N3971), .B(N5144), .CI(N4864));
ADDFX1 inst_cellmath__24_0_I1745 (.CO(N4209), .S(N3764), .A(N3088), .B(N4253), .CI(N3994));
ADDFX1 inst_cellmath__24_0_I1746 (.CO(N5112), .S(N4663), .A(N4289), .B(N4896), .CI(N3122));
ADDFX1 inst_cellmath__24_0_I1747 (.CO(N3950), .S(N3503), .A(N4929), .B(N4030), .CI(N3730));
ADDFX1 inst_cellmath__24_0_I1748 (.CO(N4849), .S(N4403), .A(N3467), .B(N4628), .CI(N3764));
ADDFX1 inst_cellmath__24_0_I1749 (.CO(N3685), .S(N3234), .A(N3503), .B(N4663), .CI(N4366));
ADDFX1 inst_cellmath__24_0_I1750 (.CO(N4589), .S(N4135), .A(N4403), .B(N3197), .CI(N4103));
ADDFX1 inst_cellmath__24_0_I1751 (.CO(N3421), .S(N5040), .A(N5006), .B(N3234), .CI(N4135));
ADDFX1 inst_cellmath__24_0_I1752 (.CO(N4321), .S(N3872), .A(N3935), .B(N4854), .CI(N4824));
ADDFX1 inst_cellmath__24_0_I1753 (.CO(N3156), .S(N4772), .A(N4549), .B(N3651), .CI(N3366));
ADDFX1 inst_cellmath__24_0_I1754 (.CO(N4060), .S(N3610), .A(N3085), .B(N4258), .CI(N3983));
ADDFX1 inst_cellmath__24_0_I1755 (.CO(N4962), .S(N4513), .A(N3697), .B(N4873), .CI(N4739));
ADDFX1 inst_cellmath__24_0_I1756 (.CO(N3800), .S(N3341), .A(N4480), .B(N3574), .CI(N3306));
ADDFX1 inst_cellmath__24_0_I1757 (.CO(N4696), .S(N4245), .A(N4772), .B(N3872), .CI(N3610));
ADDFX1 inst_cellmath__24_0_I1758 (.CO(N3534), .S(N3081), .A(N4513), .B(N4209), .CI(N5112));
ADDFX1 inst_cellmath__24_0_I1759 (.CO(N4439), .S(N3986), .A(N3950), .B(N3341), .CI(N4245));
ADDFX1 inst_cellmath__24_0_I1760 (.CO(N3264), .S(N4884), .A(N3081), .B(N4849), .CI(N3685));
ADDFX1 inst_cellmath__24_0_I1761 (.CO(N4167), .S(N3722), .A(N4589), .B(N3986), .CI(N4884));
ADDFX1 inst_cellmath__24_0_I1762 (.CO(N5074), .S(N4620), .A(N3662), .B(N3689), .CI(N4557));
ADDFX1 inst_cellmath__24_0_I1763 (.CO(N3903), .S(N3456), .A(N4267), .B(N3375), .CI(N3094));
ADDFX1 inst_cellmath__24_0_I1764 (.CO(N4806), .S(N4356), .A(N4883), .B(N3992), .CI(N3707));
ADDFX1 inst_cellmath__24_0_I1765 (.CO(N3643), .S(N3189), .A(N4321), .B(N4598), .CI(N3156));
ADDFX1 inst_cellmath__24_0_I1766 (.CO(N4547), .S(N4095), .A(N4620), .B(N4060), .CI(N3456));
ADDFX1 inst_cellmath__24_0_I1767 (.CO(N3377), .S(N4998), .A(N4962), .B(N4356), .CI(N3800));
ADDFX1 inst_cellmath__24_0_I1768 (.CO(N4280), .S(N3830), .A(N4696), .B(N3189), .CI(N4095));
ADDFX1 inst_cellmath__24_0_I1769 (.CO(N3114), .S(N4728), .A(N4998), .B(N3534), .CI(N4439));
ADDFX1 inst_cellmath__24_0_I1770 (.CO(N4019), .S(N3565), .A(N3264), .B(N3830), .CI(N4728));
ADDFX1 inst_cellmath__24_0_I1771 (.CO(N4920), .S(N4469), .A(N3387), .B(N4590), .CI(N4278));
ADDFX1 inst_cellmath__24_0_I1772 (.CO(N3755), .S(N3295), .A(N4001), .B(N3103), .CI(N4893));
ADDFX1 inst_cellmath__24_0_I1773 (.CO(N4653), .S(N4201), .A(N4607), .B(N3716), .CI(N3433));
ADDFX1 inst_cellmath__24_0_I1774 (.CO(N3493), .S(N5105), .A(N3903), .B(N5074), .CI(N4806));
ADDFX1 inst_cellmath__24_0_I1775 (.CO(N4393), .S(N3940), .A(N3295), .B(N4469), .CI(N4201));
ADDFX1 inst_cellmath__24_0_I1776 (.CO(N3225), .S(N4841), .A(N4547), .B(N3643), .CI(N5105));
ADDFX1 inst_cellmath__24_0_I1777 (.CO(N4128), .S(N3678), .A(N3940), .B(N3377), .CI(N4280));
ADDFX1 inst_cellmath__24_0_I1778 (.CO(N5033), .S(N4578), .A(N3114), .B(N4841), .CI(N3678));
ADDFX1 inst_cellmath__24_0_I1779 (.CO(N3862), .S(N3412), .A(N3116), .B(N3425), .CI(N4012));
ADDFX1 inst_cellmath__24_0_I1780 (.CO(N4763), .S(N4313), .A(N3727), .B(N4901), .CI(N4618));
ADDFX1 inst_cellmath__24_0_I1781 (.CO(N3599), .S(N3147), .A(N4332), .B(N3443), .CI(N4920));
ADDFX1 inst_cellmath__24_0_I1782 (.CO(N4503), .S(N4054), .A(N4653), .B(N3755), .CI(N3412));
ADDFX1 inst_cellmath__24_0_I1783 (.CO(N3332), .S(N4952), .A(N3493), .B(N4313), .CI(N3147));
ADDFX1 inst_cellmath__24_0_I1784 (.CO(N4236), .S(N3790), .A(N4054), .B(N4393), .CI(N3225));
ADDFX1 inst_cellmath__24_0_I1785 (.CO(N5139), .S(N4688), .A(N4128), .B(N4952), .CI(N3790));
ADDFX1 inst_cellmath__24_0_I1786 (.CO(N3976), .S(N3526), .A(N4909), .B(N4326), .CI(N3735));
ADDFX1 inst_cellmath__24_0_I1787 (.CO(N4876), .S(N4427), .A(N3453), .B(N4626), .CI(N4340));
ADDFX1 inst_cellmath__24_0_I1788 (.CO(N3712), .S(N3256), .A(N3862), .B(N3165), .CI(N4763));
ADDFX1 inst_cellmath__24_0_I1789 (.CO(N4611), .S(N4158), .A(N4427), .B(N3526), .CI(N3599));
ADDFX1 inst_cellmath__24_0_I1790 (.CO(N3446), .S(N5066), .A(N3256), .B(N4503), .CI(N3332));
ADDFX1 inst_cellmath__24_0_I1791 (.CO(N4346), .S(N3895), .A(N4236), .B(N4158), .CI(N5066));
ADDFX1 inst_cellmath__24_0_I1792 (.CO(N3181), .S(N4795), .A(N4635), .B(N3157), .CI(N3464));
ADDFX1 inst_cellmath__24_0_I1793 (.CO(N4084), .S(N3635), .A(N3178), .B(N4351), .CI(N4072));
ADDFX1 inst_cellmath__24_0_I1794 (.CO(N4991), .S(N4538), .A(N4876), .B(N3976), .CI(N4795));
ADDFX1 inst_cellmath__24_0_I1795 (.CO(N3822), .S(N3364), .A(N3712), .B(N3635), .CI(N4611));
ADDFX1 inst_cellmath__24_0_I1796 (.CO(N4720), .S(N4270), .A(N3446), .B(N4538), .CI(N3364));
ADDFX1 inst_cellmath__24_0_I1797 (.CO(N3557), .S(N3106), .A(N4362), .B(N4063), .CI(N3187));
ADDFX1 inst_cellmath__24_0_I1798 (.CO(N4461), .S(N4010), .A(N4977), .B(N4081), .CI(N3181));
ADDFX1 inst_cellmath__24_0_I1799 (.CO(N3285), .S(N4912), .A(N3106), .B(N4084), .CI(N4991));
ADDFX1 inst_cellmath__24_0_I1800 (.CO(N4193), .S(N3746), .A(N3822), .B(N4010), .CI(N4912));
ADDFX1 inst_cellmath__24_0_I1801 (.CO(N5097), .S(N4643), .A(N4090), .B(N4967), .CI(N4984));
ADDFX1 inst_cellmath__24_0_I1802 (.CO(N3932), .S(N3483), .A(N3557), .B(N3808), .CI(N4643));
ADDFX1 inst_cellmath__24_0_I1803 (.CO(N4832), .S(N4382), .A(N3483), .B(N4461), .CI(N3285));
ADDFX1 inst_cellmath__24_0_I1804 (.CO(N3670), .S(N3215), .A(N3818), .B(N3801), .CI(N4708));
ADDFX1 inst_cellmath__24_0_I1805 (.CO(N4571), .S(N4119), .A(N3215), .B(N5097), .CI(N3932));
ADDFX1 inst_cellmath__24_0_I1806 (.CO(N3690), .S(N5023), .A(N3544), .B(N4700), .CI(N3670));
NAND2XL inst_cellmath__24_0_I1807 (.Y(N3854), .A(N4178), .B(N5077));
NOR2XL inst_cellmath__24_0_I1808 (.Y(N4303), .A(N4798), .B(N4440));
NAND2XL inst_cellmath__24_0_I1809 (.Y(N4754), .A(N4798), .B(N4440));
NOR2XL inst_cellmath__24_0_I1810 (.Y(N3139), .A(N3268), .B(N4171));
NAND2XL inst_cellmath__24_0_I1811 (.Y(N3589), .A(N3268), .B(N4171));
NOR2XL inst_cellmath__24_0_I1812 (.Y(N4045), .A(N4624), .B(N4809));
NAND2XL inst_cellmath__24_0_I1813 (.Y(N4495), .A(N4624), .B(N4809));
NOR2XL inst_cellmath__24_0_I1814 (.Y(N4943), .A(N3380), .B(N4282));
NAND2X1 inst_cellmath__24_0_I1815 (.Y(N3320), .A(N3380), .B(N4282));
NOR2XL inst_cellmath__24_0_I1816 (.Y(N3782), .A(N4730), .B(N4654));
NAND2XL inst_cellmath__24_0_I1817 (.Y(N4224), .A(N4730), .B(N4654));
NOR2XL inst_cellmath__24_0_I1818 (.Y(N4678), .A(N5108), .B(N3863));
NAND2XL inst_cellmath__24_0_I1819 (.Y(N5129), .A(N5108), .B(N3863));
NOR2XL inst_cellmath__24_0_I1820 (.Y(N3517), .A(N4317), .B(N3981));
NAND2XL inst_cellmath__24_0_I1821 (.Y(N3965), .A(N4317), .B(N3981));
NOR2XL inst_cellmath__24_0_I1822 (.Y(N4418), .A(N4428), .B(N4992));
NAND2X1 inst_cellmath__24_0_I1823 (.Y(N4865), .A(N4428), .B(N4992));
NOR2X2 inst_cellmath__24_0_I1824 (.Y(N3247), .A(N3369), .B(N4834));
NAND2X1 inst_cellmath__24_0_I1825 (.Y(N3701), .A(N3369), .B(N4834));
NOR2X1 inst_cellmath__24_0_I1826 (.Y(N4148), .A(N3218), .B(N3522));
NAND2X2 inst_cellmath__24_0_I1827 (.Y(N4602), .A(N3218), .B(N3522));
NOR2XL inst_cellmath__24_0_I1828 (.Y(N5056), .A(N3970), .B(N3099));
NAND2XL inst_cellmath__24_0_I1829 (.Y(N3436), .A(N3970), .B(N3099));
NOR2X1 inst_cellmath__24_0_I1830 (.Y(N3887), .A(N3548), .B(N3585));
NAND2XL inst_cellmath__24_0_I1831 (.Y(N4336), .A(N3548), .B(N3585));
AOI21XL inst_cellmath__24_0_I1834 (.Y(N4528), .A0(N4754), .A1(N3854), .B0(N4303));
INVXL inst_cellmath__24_0_I1835 (.Y(N4226), .A(N3139));
INVXL inst_cellmath__24_0_I1836 (.Y(N4680), .A(N3589));
OAI21XL inst_cellmath__24_0_I1837 (.Y(N3999), .A0(N4680), .A1(N4528), .B0(N4226));
AOI21XL inst_cellmath__24_0_I1838 (.Y(N3473), .A0(N4495), .A1(N3999), .B0(N4045));
INVXL inst_cellmath__24_0_I1839 (.Y(N3249), .A(N4943));
INVXL inst_cellmath__24_0_I1840 (.Y(N3700), .A(N3320));
OAI21X1 inst_cellmath__24_0_I1841 (.Y(N4746), .A0(N3700), .A1(N3473), .B0(N3249));
AOI21X2 inst_cellmath__24_0_I1842 (.Y(N3954), .A0(N4224), .A1(N4746), .B0(N3782));
INVXL inst_cellmath__24_0_I1843 (.Y(N4075), .A(N4678));
INVXL inst_cellmath__24_0_I1844 (.Y(N4530), .A(N5129));
OAI21X2 inst_cellmath__24_0_I1845 (.Y(N4971), .A0(N3954), .A1(N4530), .B0(N4075));
AO21XL inst_cellmath__24_0_I1846 (.Y(N3279), .A0(N4865), .A1(N3517), .B0(N4418));
CLKAND2X2 inst_cellmath__24_0_I1847 (.Y(N3737), .A(N3965), .B(N4865));
AOI21XL inst_cellmath__24_0_I1848 (.Y(N3385), .A0(N3965), .A1(N4971), .B0(N3517));
AOI21X2 inst_cellmath__24_0_I1849 (.Y(N4286), .A0(N4971), .A1(N3737), .B0(N3279));
AOI21X2 inst_cellmath__24_0_I1850 (.Y(N4027), .A0(N4602), .A1(N3247), .B0(N4148));
NAND2X2 inst_cellmath__24_0_I1851 (.Y(N4477), .A(N4602), .B(N3701));
OAI21X2 inst_cellmath__24_0_I1852 (.Y(N3606), .A0(N4477), .A1(N4286), .B0(N4027));
NOR2BX1 inst_cellmath__24_0_I1853 (.Y(N4874), .AN(N3701), .B(N4286));
NOR2XL inst_cellmath__24_0_I1854 (.Y(N4857), .A(N4874), .B(N3247));
NAND2BXL inst_cellmath__24_0_I1862 (.Y(N5136), .AN(N4303), .B(N4754));
NAND2BXL inst_cellmath__24_0_I1863 (.Y(N4423), .AN(N3139), .B(N3589));
NAND2BXL inst_cellmath__24_0_I1864 (.Y(N3708), .AN(N4045), .B(N4495));
NAND2BXL inst_cellmath__24_0_I1865 (.Y(N5062), .AN(N4943), .B(N3320));
NAND2BXL inst_cellmath__24_0_I1866 (.Y(N4341), .AN(N3782), .B(N4224));
NAND2BXL inst_cellmath__24_0_I1867 (.Y(N3630), .AN(N4678), .B(N5129));
NAND2BXL inst_cellmath__24_0_I1868 (.Y(N4985), .AN(N3517), .B(N3965));
NAND2BXL inst_cellmath__24_0_I1869 (.Y(N4264), .AN(N4418), .B(N4865));
NAND2BXL inst_cellmath__24_0_I1870 (.Y(N3551), .AN(N3247), .B(N3701));
NAND2BXL inst_cellmath__24_0_I1871 (.Y(N4906), .AN(N4148), .B(N4602));
NAND2BXL inst_cellmath__24_0_I1872 (.Y(N4187), .AN(N5056), .B(N3436));
NAND2BXL inst_cellmath__24_0_I1873 (.Y(N3479), .AN(N3887), .B(N4336));
XNOR2X1 inst_cellmath__24_0_I1875 (.Y(inst_cellmath__24[1]), .A(N5077), .B(N4178));
XNOR2X1 inst_cellmath__24_0_I1876 (.Y(inst_cellmath__24[2]), .A(N3854), .B(N5136));
XOR2XL inst_cellmath__24_0_I1877 (.Y(inst_cellmath__24[3]), .A(N4528), .B(N4423));
XNOR2X1 inst_cellmath__24_0_I1878 (.Y(inst_cellmath__24[4]), .A(N3999), .B(N3708));
XOR2XL inst_cellmath__24_0_I1879 (.Y(inst_cellmath__24[5]), .A(N3473), .B(N5062));
XNOR2X1 inst_cellmath__24_0_I1880 (.Y(inst_cellmath__24[6]), .A(N4746), .B(N4341));
XOR2XL inst_cellmath__24_0_I1881 (.Y(inst_cellmath__24[7]), .A(N3954), .B(N3630));
XNOR2X1 inst_cellmath__24_0_I1882 (.Y(inst_cellmath__24[8]), .A(N4971), .B(N4985));
CLKXOR2X1 inst_cellmath__24_0_I1883 (.Y(inst_cellmath__24[9]), .A(N3385), .B(N4264));
XOR2XL inst_cellmath__24_0_I1884 (.Y(inst_cellmath__24[10]), .A(N4286), .B(N3551));
XOR2XL inst_cellmath__24_0_I1885 (.Y(inst_cellmath__24[11]), .A(N4857), .B(N4906));
XNOR2X1 inst_cellmath__24_0_I1886 (.Y(inst_cellmath__24[12]), .A(N3606), .B(N4187));
AOI21X2 inst_cellmath__25_0_I13760 (.Y(N4092), .A0(N3436), .A1(N3606), .B0(N5056));
XOR2XL inst_cellmath__24_0_I1887 (.Y(inst_cellmath__24[13]), .A(N4092), .B(N3479));
NOR2X2 inst_cellmath__24_0_I1891 (.Y(N3514), .A(N3575), .B(N4246));
NAND2X1 inst_cellmath__24_0_I1892 (.Y(N3962), .A(N3575), .B(N4246));
NOR2X1 inst_cellmath__24_0_I1893 (.Y(N4415), .A(N4697), .B(N4202));
NAND2X2 inst_cellmath__24_0_I1894 (.Y(N4862), .A(N4697), .B(N4202));
NOR2X1 inst_cellmath__24_0_I1895 (.Y(N3243), .A(N4652), .B(N5064));
NAND2X2 inst_cellmath__24_0_I1896 (.Y(N3698), .A(N4652), .B(N5064));
NOR2XL inst_cellmath__24_0_I1897 (.Y(N4146), .A(N3447), .B(N4755));
NAND2X4 inst_cellmath__24_0_I1898 (.Y(N4599), .A(N3447), .B(N4755));
NAND2XL inst_cellmath__24_0_I1900 (.Y(N3431), .A(N3136), .B(N3278));
ADDFHXL inst_cellmath__24_0_I13824 (.CO(N4725), .S(N22739), .A(N4658), .B(N4546), .CI(N3370));
NOR2X2 inst_cellmath__24_0_I1907 (.Y(N4524), .A(N4725), .B(N3442));
NAND2XL inst_cellmath__24_0_I1908 (.Y(N4978), .A(N4725), .B(N3442));
NOR2X1 inst_cellmath__24_0_I1909 (.Y(N3353), .A(N3892), .B(N3777));
NAND2X2 inst_cellmath__24_0_I1910 (.Y(N3809), .A(N3892), .B(N3777));
NOR2X2 inst_cellmath__24_0_I1911 (.Y(N4256), .A(N4221), .B(N3200));
NAND2X2 inst_cellmath__24_0_I1912 (.Y(N4706), .A(N4221), .B(N3200));
NOR2XL inst_cellmath__24_0_I1913 (.Y(N3092), .A(N3658), .B(N3802));
NAND2X2 inst_cellmath__24_0_I1914 (.Y(N3545), .A(N3658), .B(N3802));
NOR2X2 inst_cellmath__24_0_I1915 (.Y(N3997), .A(N4247), .B(N3498));
NAND2X1 inst_cellmath__24_0_I1916 (.Y(N4449), .A(N4247), .B(N3498));
NOR2X1 inst_cellmath__24_0_I1917 (.Y(N4899), .A(N3943), .B(N4350));
NAND2X2 inst_cellmath__24_0_I1918 (.Y(N3275), .A(N3943), .B(N4350));
NOR2X1 inst_cellmath__24_0_I1919 (.Y(N3733), .A(N4799), .B(N4307));
NAND2X2 inst_cellmath__24_0_I1920 (.Y(N4179), .A(N4799), .B(N4307));
NOR2XL inst_cellmath__24_0_I1921 (.Y(N4631), .A(N4759), .B(N3359));
NAND2X2 inst_cellmath__24_0_I1922 (.Y(N5085), .A(N4759), .B(N3359));
NOR2X2 inst_cellmath__24_0_I1923 (.Y(N3470), .A(N3815), .B(N3584));
NAND2X1 inst_cellmath__24_0_I1924 (.Y(N3919), .A(N3815), .B(N3584));
NOR2X1 inst_cellmath__24_0_I1925 (.Y(N4369), .A(N4039), .B(N4974));
NAND2X2 inst_cellmath__24_0_I1926 (.Y(N4818), .A(N4039), .B(N4974));
NOR2X1 inst_cellmath__24_0_I1927 (.Y(N3203), .A(N3350), .B(N3388));
NAND2X1 inst_cellmath__24_0_I1928 (.Y(N3657), .A(N3350), .B(N3388));
NOR2XL inst_cellmath__24_0_I1929 (.Y(N4106), .A(N3839), .B(N5040));
NAND2X2 inst_cellmath__24_0_I1930 (.Y(N4560), .A(N3839), .B(N5040));
NOR2XL inst_cellmath__24_0_I1931 (.Y(N5010), .A(N3421), .B(N3722));
NAND2XL inst_cellmath__24_0_I1932 (.Y(N3391), .A(N3421), .B(N3722));
NOR2XL inst_cellmath__24_0_I1933 (.Y(N3844), .A(N4167), .B(N3565));
NAND2XL inst_cellmath__24_0_I1934 (.Y(N4293), .A(N4167), .B(N3565));
NOR2XL inst_cellmath__24_0_I1935 (.Y(N4742), .A(N4019), .B(N4578));
NAND2XL inst_cellmath__24_0_I1936 (.Y(N3126), .A(N4019), .B(N4578));
NOR2XL inst_cellmath__24_0_I1937 (.Y(N3577), .A(N5033), .B(N4688));
NAND2XL inst_cellmath__24_0_I1938 (.Y(N4032), .A(N5033), .B(N4688));
NOR2XL inst_cellmath__24_0_I1939 (.Y(N4485), .A(N5139), .B(N3895));
NAND2XL inst_cellmath__24_0_I1940 (.Y(N4933), .A(N5139), .B(N3895));
NOR2XL inst_cellmath__24_0_I1941 (.Y(N3308), .A(N4346), .B(N4270));
NAND2XL inst_cellmath__24_0_I1942 (.Y(N3770), .A(N4346), .B(N4270));
NOR2XL inst_cellmath__24_0_I1943 (.Y(N4211), .A(N4720), .B(N3746));
NAND2XL inst_cellmath__24_0_I1944 (.Y(N4665), .A(N4720), .B(N3746));
NOR2XL inst_cellmath__24_0_I1945 (.Y(N5117), .A(N4382), .B(N4193));
NAND2XL inst_cellmath__24_0_I1946 (.Y(N3506), .A(N4382), .B(N4193));
NOR2XL inst_cellmath__24_0_I1947 (.Y(N3952), .A(N4119), .B(N4832));
NAND2XL inst_cellmath__24_0_I1948 (.Y(N4407), .A(N4119), .B(N4832));
NOR2XL inst_cellmath__24_0_I1949 (.Y(N4852), .A(N5023), .B(N4571));
NAND2XL inst_cellmath__24_0_I1950 (.Y(N3236), .A(N5023), .B(N4571));
NAND2X1 inst_cellmath__25_0_I13771 (.Y(N5126), .A(N3351), .B(N3123));
NAND2X2 inst_cellmath__25_0_I13759 (.Y(N22575), .A(N4038), .B(N4972));
NAND2X1 inst_cellmath__25_0_I13763 (.Y(N22578), .A(N4336), .B(N22575));
NOR2XL inst_cellmath__25_0_I13758 (.Y(N22566), .A(N4038), .B(N4972));
AOI21X1 inst_cellmath__25_0_I13762 (.Y(N22570), .A0(N3887), .A1(N22575), .B0(N22566));
OAI21X2 inst_cellmath__25_0_I13766 (.Y(N3778), .A0(N22578), .A1(N4092), .B0(N22570));
NOR2XL inst_cellmath__25_0_I13770 (.Y(N4674), .A(N3351), .B(N3123));
AOI21X2 inst_cellmath__24_0_I1951 (.Y(N5045), .A0(N5126), .A1(N3778), .B0(N4674));
AOI21X2 inst_cellmath__24_0_I1952 (.Y(N4776), .A0(N3514), .A1(N4862), .B0(N4415));
NAND2X2 inst_cellmath__24_0_I1953 (.Y(N3158), .A(N3962), .B(N4862));
INVXL inst_cellmath__24_0_I1954 (.Y(N3618), .A(N3243));
INVXL inst_cellmath__24_0_I1955 (.Y(N4066), .A(N3698));
AOI21X2 inst_cellmath__24_0_I1956 (.Y(N4516), .A0(N3243), .A1(N4599), .B0(N4146));
NAND2X4 inst_cellmath__24_0_I1957 (.Y(N4968), .A(N3698), .B(N4599));
INVXL inst_cellmath__24_0_I1958 (.Y(N3349), .A(N4776));
OAI21XL inst_cellmath__24_0_I1959 (.Y(N3083), .A0(N4066), .A1(N4776), .B0(N3618));
AOI21X2 inst_cellmath__24_0_I1965 (.Y(N3192), .A0(N3809), .A1(N4524), .B0(N3353));
AOI21X1 inst_cellmath__24_0_I1966 (.Y(N5002), .A0(N4256), .A1(N3545), .B0(N3092));
AOI21X2 inst_cellmath__24_0_I1968 (.Y(N4732), .A0(N3997), .A1(N3275), .B0(N4899));
AOI21XL inst_cellmath__24_0_I1969 (.Y(N4473), .A0(N5085), .A1(N3733), .B0(N4631));
AOI21X2 inst_cellmath__24_0_I1970 (.Y(N4204), .A0(N4818), .A1(N3470), .B0(N4369));
NAND2X1 inst_cellmath__24_0_I1971 (.Y(N4656), .A(N4818), .B(N3919));
INVXL inst_cellmath__24_0_I1972 (.Y(N4364), .A(N3203));
INVXL inst_cellmath__24_0_I1973 (.Y(N4812), .A(N3657));
AOI21X1 inst_cellmath__24_0_I1974 (.Y(N3942), .A0(N3203), .A1(N4560), .B0(N4106));
NAND2X2 inst_cellmath__24_0_I1975 (.Y(N4399), .A(N4560), .B(N3657));
INVXL inst_cellmath__24_0_I1976 (.Y(N4100), .A(N4204));
OAI21XL inst_cellmath__24_0_I1977 (.Y(N4580), .A0(N4812), .A1(N4204), .B0(N4364));
OAI21X4 inst_cellmath__24_0_I1978 (.Y(N3414), .A0(N4399), .A1(N4204), .B0(N3942));
NOR2X1 inst_cellmath__24_0_I1979 (.Y(N3866), .A(N4399), .B(N4656));
AOI21X1 inst_cellmath__24_0_I1980 (.Y(N3149), .A0(N4293), .A1(N5010), .B0(N3844));
NAND2X1 inst_cellmath__24_0_I1981 (.Y(N3605), .A(N4293), .B(N3391));
INVXL inst_cellmath__24_0_I1982 (.Y(N3837), .A(N4742));
INVXL inst_cellmath__24_0_I1983 (.Y(N4288), .A(N3126));
AOI21XL inst_cellmath__24_0_I1984 (.Y(N4958), .A0(N4032), .A1(N4742), .B0(N3577));
NAND2XL inst_cellmath__24_0_I1985 (.Y(N3336), .A(N4032), .B(N3126));
INVXL inst_cellmath__24_0_I1986 (.Y(N3572), .A(N3149));
OAI21XL inst_cellmath__24_0_I1987 (.Y(N3531), .A0(N4288), .A1(N3149), .B0(N3837));
OAI21X1 inst_cellmath__24_0_I1988 (.Y(N4430), .A0(N3336), .A1(N3149), .B0(N4958));
NOR2X1 inst_cellmath__24_0_I1989 (.Y(N4881), .A(N3336), .B(N3605));
AOI21XL inst_cellmath__24_0_I1990 (.Y(N4163), .A0(N3770), .A1(N4485), .B0(N3308));
NAND2XL inst_cellmath__24_0_I1991 (.Y(N4614), .A(N3770), .B(N4933));
INVXL inst_cellmath__24_0_I1992 (.Y(N3301), .A(N4211));
INVXL inst_cellmath__24_0_I1993 (.Y(N3763), .A(N4665));
AOI21XL inst_cellmath__24_0_I1994 (.Y(N3897), .A0(N3506), .A1(N4211), .B0(N5117));
NAND2XL inst_cellmath__24_0_I1995 (.Y(N4349), .A(N3506), .B(N4665));
INVXL inst_cellmath__24_0_I1996 (.Y(N5110), .A(N4163));
OAI21XL inst_cellmath__24_0_I1997 (.Y(N4542), .A0(N3763), .A1(N4163), .B0(N3301));
AOI21XL inst_cellmath__24_0_I1998 (.Y(N3109), .A0(N3236), .A1(N3952), .B0(N4852));
NAND2XL inst_cellmath__24_0_I1999 (.Y(N3560), .A(N3236), .B(N4407));
INVXL inst_cellmath__24_0_I2000 (.Y(N4584), .A(N3109));
NOR2X2 inst_cellmath__24_0_I2001 (.Y(N4002), .A(N3690), .B(N3109));
NOR2X1 inst_cellmath__24_0_I2002 (.Y(N3487), .A(N3690), .B(N3560));
ADDFHX1 inst_cellmath__24_0_I13822 (.CO(N22749), .S(N22743), .A(N4900), .B(N5046), .CI(N3877));
NAND2X2 inst_cellmath__24_0_I13827 (.Y(N4333), .A(N3736), .B(N22743));
INVX2 inst_cellmath__24_0_I13929 (.Y(N3418), .A(N5045));
INVXL inst_cellmath__24_0_I2016 (.Y(N4353), .A(N3418));
CLKAND2X2 inst_cellmath__24_0_I13930 (.Y(N3151), .A(N3431), .B(N4333));
INVXL inst_cellmath__24_0_I2018 (.Y(N4091), .A(N3151));
ADDFHXL inst_cellmath__24_0_I13823 (.CO(N22731), .S(N22757), .A(N4327), .B(N3300), .CI(N4207));
NOR2X2 inst_cellmath__24_0_I13825 (.Y(N5053), .A(N3136), .B(N3278));
NOR2X1 inst_cellmath__24_0_I13826 (.Y(N3883), .A(N3736), .B(N22743));
NOR2X2 inst_cellmath__24_0_I13828 (.Y(N4783), .A(N22749), .B(N22757));
NAND2X2 inst_cellmath__24_0_I13829 (.Y(N3166), .A(N22749), .B(N22757));
NOR2XL inst_cellmath__24_0_I13830 (.Y(N3624), .A(N22731), .B(N22739));
NAND2X2 inst_cellmath__24_0_I13831 (.Y(N22759), .A(N22731), .B(N22739));
AOI21X2 inst_cellmath__24_0_I13832 (.Y(N22737), .A0(N5053), .A1(N4333), .B0(N3883));
AOI21X2 inst_cellmath__24_0_I13833 (.Y(N22745), .A0(N4783), .A1(N22759), .B0(N3624));
OAI21X2 inst_cellmath__24_0_I13926 (.Y(N22911), .A0(N4968), .A1(N4776), .B0(N4516));
NOR2X2 inst_cellmath__24_0_I13927 (.Y(N22921), .A(N3158), .B(N4968));
CLKAND2X3 inst_cellmath__24_0_I13928 (.Y(N22933), .A(N3545), .B(N4706));
CLKINVX2 inst_cellmath__24_0_I13931 (.Y(N4244), .A(N3192));
CLKAND2X2 inst_cellmath__24_0_I13932 (.Y(N4694), .A(N4978), .B(N3809));
CLKINVX1 inst_cellmath__24_0_I13933 (.Y(N22938), .A(N5002));
INVX2 inst_cellmath__24_0_I13934 (.Y(N3718), .A(N4732));
CLKAND2X3 inst_cellmath__24_0_I13935 (.Y(N4166), .A(N3275), .B(N4449));
INVX1 inst_cellmath__24_0_I13936 (.Y(N22919), .A(N4473));
CLKAND2X3 inst_cellmath__24_0_I13937 (.Y(N22931), .A(N5085), .B(N4179));
AOI21X4 inst_cellmath__24_0_I13938 (.Y(N5058), .A0(N22921), .A1(N3418), .B0(N22911));
CLKAND2X6 inst_cellmath__24_0_I13939 (.Y(N22951), .A(N3166), .B(N22759));
NAND2X4 inst_cellmath__24_0_I13940 (.Y(N22954), .A(N3151), .B(N22951));
INVX2 inst_cellmath__24_0_I13941 (.Y(N4771), .A(N22737));
INVX2 inst_cellmath__24_0_I13942 (.Y(N22922), .A(N22745));
AOI21X4 inst_cellmath__24_0_I13943 (.Y(N22934), .A0(N4771), .A1(N22951), .B0(N22922));
OAI21X4 inst_cellmath__24_0_I13944 (.Y(N4261), .A0(N22954), .A1(N5058), .B0(N22934));
AOI21X4 inst_cellmath__24_0_I13945 (.Y(N22915), .A0(N22933), .A1(N4244), .B0(N22938));
NAND2X4 inst_cellmath__24_0_I13946 (.Y(N4454), .A(N4694), .B(N22933));
AOI21X4 inst_cellmath__24_0_I13947 (.Y(N22947), .A0(N22931), .A1(N3718), .B0(N22919));
NAND2X6 inst_cellmath__24_0_I13948 (.Y(N22958), .A(N22931), .B(N4166));
OAI21X4 inst_cellmath__24_0_I13949 (.Y(N22917), .A0(N22958), .A1(N22915), .B0(N22947));
NOR2X4 inst_cellmath__24_0_I13950 (.Y(N22928), .A(N22958), .B(N4454));
AOI21X4 inst_cellmath__24_0_I13951 (.Y(N4218), .A0(N4261), .A1(N22928), .B0(N22917));
DLY1X1 inst_cellmath__24_0_I13952 (.Y(N4006), .A(N22915));
INVXL inst_cellmath__24_0_I2024 (.Y(N4918), .A(N3718));
INVXL inst_cellmath__24_0_I2025 (.Y(N3292), .A(N4166));
INVXL inst_cellmath__24_0_I2028 (.Y(N4651), .A(N4006));
INVXL inst_cellmath__24_0_I2029 (.Y(N5103), .A(N4454));
OAI21X1 inst_cellmath__24_0_I2030 (.Y(N4375), .A0(N3292), .A1(N4006), .B0(N4918));
NOR2XL inst_cellmath__24_0_I2031 (.Y(N4825), .A(N3292), .B(N4454));
NOR2XL inst_cellmath__24_0_I2034 (.Y(N3434), .A(N4091), .B(N5058));
NOR2XL inst_cellmath__24_0_I2035 (.Y(N4392), .A(N3434), .B(N4771));
INVXL buf1_A_I5419 (.Y(N11836), .A(N4261));
INVXL buf1_A_I5420 (.Y(N4837), .A(N11836));
AOI21XL inst_cellmath__24_0_I2037 (.Y(N3583), .A0(N4694), .A1(N4261), .B0(N4244));
AOI21XL inst_cellmath__24_0_I2038 (.Y(N4491), .A0(N5103), .A1(N4261), .B0(N4651));
AOI21XL inst_cellmath__24_0_I2039 (.Y(N3315), .A0(N4825), .A1(N4261), .B0(N4375));
AOI21X4 inst_cellmath__24_0_I2043 (.Y(N3959), .A0(N4881), .A1(N3414), .B0(N4430));
NAND2XL inst_cellmath__24_0_I2044 (.Y(N4412), .A(N4881), .B(N3866));
OA21X1 inst_cellmath__24_0_I2045 (.Y(N5032), .A0(N4349), .A1(N4163), .B0(N3897));
OR2XL inst_cellmath__24_0_I2046 (.Y(N3408), .A(N4349), .B(N4614));
OAI21X2 inst_cellmath__24_0_I2047 (.Y(N3427), .A0(N3408), .A1(N3959), .B0(N5032));
INVXL inst_cellmath__24_0_I2048 (.Y(N3598), .A(N3414));
INVXL inst_cellmath__24_0_I2049 (.Y(N4050), .A(N3866));
INVX2 inst_cellmath__24_0_I2050 (.Y(N3328), .A(N3427));
OR2X1 inst_cellmath__24_0_I2051 (.Y(N3786), .A(N3408), .B(N4412));
OAI21XL inst_cellmath__24_0_I2052 (.Y(N3916), .A0(N4050), .A1(N4218), .B0(N3598));
OAI21X4 inst_cellmath__24_0_I2054 (.Y(N3652), .A0(N3786), .A1(N4218), .B0(N3328));
NAND2BXL inst_cellmath__24_0_I2057 (.Y(N4029), .AN(N3514), .B(N3962));
NAND2BXL inst_cellmath__24_0_I2058 (.Y(N3305), .AN(N4415), .B(N4862));
NAND2BXL inst_cellmath__24_0_I2059 (.Y(N4662), .AN(N3243), .B(N3698));
NAND2BXL inst_cellmath__24_0_I2060 (.Y(N3949), .AN(N4146), .B(N4599));
NAND2BXL inst_cellmath__24_0_I2061 (.Y(N3233), .AN(N5053), .B(N3431));
NAND2BXL inst_cellmath__24_0_I2062 (.Y(N4588), .AN(N3883), .B(N4333));
NAND2BXL inst_cellmath__24_0_I2063 (.Y(N3871), .AN(N4783), .B(N3166));
NAND2BXL inst_cellmath__24_0_I13980 (.Y(N3155), .AN(N3624), .B(N22759));
NAND2BXL inst_cellmath__24_0_I2065 (.Y(N4512), .AN(N4524), .B(N4978));
NAND2BXL inst_cellmath__24_0_I2066 (.Y(N3799), .AN(N3353), .B(N3809));
NAND2BXL inst_cellmath__24_0_I2067 (.Y(N3080), .AN(N4256), .B(N4706));
NAND2BXL inst_cellmath__24_0_I2068 (.Y(N4438), .AN(N3092), .B(N3545));
NAND2BXL inst_cellmath__24_0_I2069 (.Y(N3721), .AN(N3997), .B(N4449));
NAND2BXL inst_cellmath__24_0_I2070 (.Y(N5073), .AN(N4899), .B(N3275));
NAND2BXL inst_cellmath__24_0_I2071 (.Y(N4355), .AN(N3733), .B(N4179));
NAND2BXL inst_cellmath__24_0_I2072 (.Y(N3642), .AN(N4631), .B(N5085));
NAND2BXL inst_cellmath__24_0_I2073 (.Y(N4997), .AN(N3470), .B(N3919));
NAND2BXL inst_cellmath__24_0_I2074 (.Y(N4279), .AN(N4369), .B(N4818));
NAND2BXL inst_cellmath__24_0_I2075 (.Y(N3564), .AN(N3203), .B(N3657));
NAND2BXL inst_cellmath__24_0_I2076 (.Y(N4919), .AN(N4106), .B(N4560));
NAND2BXL inst_cellmath__24_0_I2077 (.Y(N4200), .AN(N5010), .B(N3391));
NAND2BXL inst_cellmath__24_0_I2078 (.Y(N3492), .AN(N3844), .B(N4293));
NAND2BXL inst_cellmath__24_0_I2079 (.Y(N4840), .AN(N4742), .B(N3126));
NAND2BXL inst_cellmath__24_0_I2080 (.Y(N4127), .AN(N3577), .B(N4032));
NAND2BXL inst_cellmath__24_0_I2081 (.Y(N3411), .AN(N4485), .B(N4933));
NAND2BXL inst_cellmath__24_0_I2082 (.Y(N4762), .AN(N3308), .B(N3770));
NAND2BXL inst_cellmath__24_0_I2083 (.Y(N4053), .AN(N4211), .B(N4665));
NAND2BXL inst_cellmath__24_0_I2084 (.Y(N3331), .AN(N5117), .B(N3506));
NAND2BXL inst_cellmath__24_0_I2086 (.Y(N3975), .AN(N4852), .B(N3236));
XOR2XL inst_cellmath__24_0_I2088 (.Y(inst_cellmath__24[16]), .A(N4353), .B(N4029));
XOR2XL inst_cellmath__24_0_I2089 (.Y(inst_cellmath__24[20]), .A(N5058), .B(N3233));
XNOR2X1 inst_cellmath__24_0_I2091 (.Y(inst_cellmath__24[24]), .A(N4837), .B(N4512));
XOR2XL inst_cellmath__24_0_I2092 (.Y(inst_cellmath__24[26]), .A(N3583), .B(N3080));
XOR2XL inst_cellmath__24_0_I2093 (.Y(inst_cellmath__24[28]), .A(N4491), .B(N3721));
XOR2XL inst_cellmath__24_0_I2094 (.Y(inst_cellmath__24[30]), .A(N3315), .B(N4355));
XOR2XL inst_cellmath__24_0_I2095 (.Y(inst_cellmath__24[32]), .A(N4218), .B(N4997));
XNOR2X1 inst_cellmath__24_0_I2096 (.Y(inst_cellmath__24[36]), .A(N4200), .B(N3916));
OAI21X1 inst_cellmath__25_0_I13875 (.Y(N4815), .A0(N4412), .A1(N4218), .B0(N3959));
XNOR2X1 inst_cellmath__24_0_I2097 (.Y(inst_cellmath__24[40]), .A(N4815), .B(N3411));
XNOR2X1 inst_cellmath__24_0_I2099 (.Y(N3821), .A(N3962), .B(N3305));
XNOR2X1 inst_cellmath__24_0_I2100 (.Y(N4269), .A(N3514), .B(N3305));
MX2XL inst_cellmath__24_0_I2101 (.Y(inst_cellmath__24[17]), .A(N3821), .B(N4269), .S0(N4353));
XNOR2X1 inst_cellmath__24_0_I2102 (.Y(N3105), .A(N4662), .B(N3349));
NOR2BX1 inst_cellmath__24_0_I2103 (.Y(N3455), .AN(N3158), .B(N3349));
XOR2XL inst_cellmath__24_0_I2104 (.Y(N3556), .A(N4662), .B(N3455));
MX2XL inst_cellmath__24_0_I2105 (.Y(inst_cellmath__24[18]), .A(N3556), .B(N3105), .S0(N4353));
XNOR2X1 inst_cellmath__24_0_I2106 (.Y(N4460), .A(N3949), .B(N3083));
NOR2XL inst_cellmath__24_0_I2107 (.Y(N5093), .A(N4066), .B(N3158));
NOR2XL inst_cellmath__24_0_I2108 (.Y(N3373), .A(N5093), .B(N3083));
XOR2XL inst_cellmath__24_0_I2109 (.Y(N4911), .A(N3949), .B(N3373));
MX2XL inst_cellmath__24_0_I2110 (.Y(inst_cellmath__24[19]), .A(N4911), .B(N4460), .S0(N4353));
XNOR2X1 inst_cellmath__24_0_I2111 (.Y(N3745), .A(N3431), .B(N4588));
XNOR2X1 inst_cellmath__24_0_I2112 (.Y(N4192), .A(N5053), .B(N4588));
MX2XL inst_cellmath__24_0_I2113 (.Y(inst_cellmath__24[21]), .A(N3745), .B(N4192), .S0(N5058));
XNOR2X1 inst_cellmath__24_0_I2114 (.Y(N5096), .A(N3166), .B(N3155));
XNOR2X1 inst_cellmath__24_0_I2115 (.Y(N3482), .A(N4783), .B(N3155));
XNOR2X1 inst_cellmath__24_0_I2117 (.Y(N4384), .A(N4978), .B(N3799));
XNOR2X1 inst_cellmath__24_0_I2118 (.Y(N4831), .A(N4524), .B(N3799));
MX2XL inst_cellmath__24_0_I2119 (.Y(inst_cellmath__24[25]), .A(N4831), .B(N4384), .S0(N4837));
XNOR2X1 inst_cellmath__24_0_I2120 (.Y(N3672), .A(N4706), .B(N4438));
XNOR2X1 inst_cellmath__24_0_I2121 (.Y(N4118), .A(N4256), .B(N4438));
MX2XL inst_cellmath__24_0_I2122 (.Y(inst_cellmath__24[27]), .A(N3672), .B(N4118), .S0(N3583));
XNOR2X1 inst_cellmath__24_0_I2123 (.Y(N5025), .A(N4449), .B(N5073));
XNOR2X1 inst_cellmath__24_0_I2124 (.Y(N3402), .A(N3997), .B(N5073));
MX2XL inst_cellmath__24_0_I2125 (.Y(inst_cellmath__24[29]), .A(N5025), .B(N3402), .S0(N4491));
XNOR2X1 inst_cellmath__24_0_I2126 (.Y(N4306), .A(N4179), .B(N3642));
XNOR2X1 inst_cellmath__24_0_I2127 (.Y(N4753), .A(N3733), .B(N3642));
MX2XL inst_cellmath__24_0_I2128 (.Y(inst_cellmath__24[31]), .A(N4306), .B(N4753), .S0(N3315));
XNOR2X1 inst_cellmath__24_0_I2129 (.Y(N3591), .A(N4279), .B(N3919));
XNOR2X1 inst_cellmath__24_0_I2130 (.Y(N4044), .A(N4279), .B(N3470));
MX2XL inst_cellmath__24_0_I2131 (.Y(inst_cellmath__24[33]), .A(N3591), .B(N4044), .S0(N4218));
XNOR2X1 inst_cellmath__24_0_I2132 (.Y(N4947), .A(N3564), .B(N4100));
NOR2BX1 inst_cellmath__24_0_I2133 (.Y(N4717), .AN(N4656), .B(N4100));
XOR2XL inst_cellmath__24_0_I2134 (.Y(N3319), .A(N3564), .B(N4717));
MX2XL inst_cellmath__24_0_I2135 (.Y(inst_cellmath__24[34]), .A(N3319), .B(N4947), .S0(N4218));
XNOR2X1 inst_cellmath__24_0_I2136 (.Y(N4227), .A(N4919), .B(N4580));
NOR2XL inst_cellmath__24_0_I2137 (.Y(N4116), .A(N4812), .B(N4656));
NOR2XL inst_cellmath__24_0_I2138 (.Y(N4641), .A(N4116), .B(N4580));
XOR2XL inst_cellmath__24_0_I2139 (.Y(N4677), .A(N4919), .B(N4641));
MX2XL inst_cellmath__24_0_I2140 (.Y(inst_cellmath__24[35]), .A(N4677), .B(N4227), .S0(N4218));
XNOR2X1 inst_cellmath__24_0_I2141 (.Y(N3520), .A(N3492), .B(N3391));
XNOR2X1 inst_cellmath__24_0_I2142 (.Y(N3964), .A(N3492), .B(N5010));
MX2XL inst_cellmath__24_0_I2143 (.Y(inst_cellmath__24[37]), .A(N3964), .B(N3520), .S0(N3916));
XNOR2X1 inst_cellmath__24_0_I2144 (.Y(N4867), .A(N4840), .B(N3572));
NOR2BX1 inst_cellmath__24_0_I2145 (.Y(N3588), .AN(N3605), .B(N3572));
XOR2XL inst_cellmath__24_0_I2146 (.Y(N3246), .A(N4840), .B(N3588));
MX2XL inst_cellmath__24_0_I2147 (.Y(inst_cellmath__24[38]), .A(N4867), .B(N3246), .S0(N3916));
XNOR2X1 inst_cellmath__24_0_I2148 (.Y(N4151), .A(N4127), .B(N3531));
NOR2XL inst_cellmath__24_0_I2149 (.Y(N3135), .A(N4288), .B(N3605));
NOR2XL inst_cellmath__24_0_I2150 (.Y(N3516), .A(N3135), .B(N3531));
XOR2XL inst_cellmath__24_0_I2151 (.Y(N4601), .A(N4127), .B(N3516));
MX2XL inst_cellmath__24_0_I2152 (.Y(inst_cellmath__24[39]), .A(N4151), .B(N4601), .S0(N3916));
XNOR2X1 inst_cellmath__24_0_I2153 (.Y(N3438), .A(N4762), .B(N4933));
XNOR2X1 inst_cellmath__24_0_I2154 (.Y(N3886), .A(N4762), .B(N4485));
MX2XL inst_cellmath__24_0_I2155 (.Y(inst_cellmath__24[41]), .A(N3886), .B(N3438), .S0(N4815));
XNOR2X1 inst_cellmath__24_0_I2156 (.Y(N4788), .A(N4053), .B(N5110));
NOR2BX1 inst_cellmath__24_0_I2157 (.Y(N4523), .AN(N4614), .B(N5110));
XOR2XL inst_cellmath__24_0_I2158 (.Y(N3169), .A(N4053), .B(N4523));
MX2XL inst_cellmath__24_0_I2159 (.Y(inst_cellmath__24[42]), .A(N4788), .B(N3169), .S0(N4815));
NOR2XL inst_cellmath__24_0_I2161 (.Y(N4223), .A(N3763), .B(N4614));
NOR2XL inst_cellmath__24_0_I2162 (.Y(N4448), .A(N4223), .B(N4542));
XNOR2X1 inst_cellmath__24_0_I2168 (.Y(N4711), .A(N3690), .B(N4584));
NOR2BX1 inst_cellmath__24_0_I2169 (.Y(N3390), .AN(N3560), .B(N4584));
XOR2XL inst_cellmath__24_0_I2170 (.Y(N3095), .A(N3690), .B(N3390));
INVXL inst_cellmath__25_0_I13876 (.Y(N3973), .A(N3652));
MX2XL inst_cellmath__24_0_I2171 (.Y(inst_cellmath__24[46]), .A(N3095), .B(N4711), .S0(N3973));
AOI21X4 inst_cellmath__25_0_I13774 (.Y(inst_cellmath__24[47]), .A0(N3487), .A1(N3652), .B0(N4002));
NAND2BXL inst_cellmath__25_0_I13877 (.Y(N22795), .AN(N3952), .B(N4407));
XNOR2X1 inst_cellmath__25_0_I13982 (.Y(N22818), .A(N22795), .B(N3973));
XOR2XL inst_cellmath__25_0_I13880 (.Y(N22802), .A(N3973), .B(N22795));
XNOR2X1 inst_cellmath__25_0_I13881 (.Y(N22810), .A(N3331), .B(N4542));
XOR2XL inst_cellmath__25_0_I13882 (.Y(N22816), .A(N3331), .B(N4448));
INVX1 inst_cellmath__25_0_I13883 (.Y(N22819), .A(N4815));
MXI2XL inst_cellmath__25_0_I13884 (.Y(N22804), .A(N22816), .B(N22810), .S0(N22819));
MX2XL inst_cellmath__25_0_I13885 (.Y(inst_cellmath__24[43]), .A(N22816), .B(N22810), .S0(N22819));
XNOR2X1 inst_cellmath__25_0_I13886 (.Y(N22798), .A(N4407), .B(N3975));
XNOR2X1 inst_cellmath__25_0_I13887 (.Y(N22806), .A(N3975), .B(N3952));
MXI2XL inst_cellmath__25_0_I13888 (.Y(N22815), .A(N22798), .B(N22806), .S0(N3973));
MX2XL inst_cellmath__25_0_I13889 (.Y(inst_cellmath__24[45]), .A(N22798), .B(N22806), .S0(N3973));
INVX6 inst_cellmath__25_0_I13890 (.Y(N11799), .A(inst_cellmath__24[47]));
INVX1 inst_cellmath__25_0_I13891 (.Y(N11806), .A(N11799));
MXI2XL inst_cellmath__25_0_I13892 (.Y(inst_cellmath__25[44]), .A(inst_cellmath__24[43]), .B(N22802), .S0(N11806));
MXI2XL inst_cellmath__25_0_I13893 (.Y(inst_cellmath__25[45]), .A(N22802), .B(inst_cellmath__24[45]), .S0(N11806));
MXI2XL inst_cellmath__25_0_I13894 (.Y(N22788), .A(N22818), .B(N22815), .S0(N11806));
MXI2XL inst_cellmath__25_0_I13895 (.Y(N22792), .A(N22804), .B(N22818), .S0(N11806));
NOR2XL inst_cellmath__25_0_I13896 (.Y(N7419), .A(N22788), .B(N22792));
INVX2 inst_cellmath__25_0_I5136 (.Y(N11807), .A(N11799));
INVXL inst_cellmath__25_0_I5133 (.Y(N11804), .A(N11799));
INVXL inst_cellmath__25_0_I5132 (.Y(N11803), .A(N11799));
CLKINVX3 inst_cellmath__25_0_I5131 (.Y(N11802), .A(N11799));
NOR2BX1 inst_cellmath__25_0_I13983 (.Y(N22579), .AN(N4336), .B(N4092));
NOR2XL inst_cellmath__25_0_I13765 (.Y(N22563), .A(N3887), .B(N22579));
NOR2BX1 inst_cellmath__25_0_I13984 (.Y(N22569), .AN(N22575), .B(N22566));
XNOR2X1 inst_cellmath__25_0_I13769 (.Y(inst_cellmath__24[14]), .A(N22569), .B(N22563));
NAND2BXL inst_cellmath__25_0_I13772 (.Y(N22560), .AN(N4674), .B(N5126));
XNOR2X1 inst_cellmath__25_0_I13773 (.Y(inst_cellmath__24[15]), .A(N3778), .B(N22560));
INVX1 inst_cellmath__25_0_I13776 (.Y(N11801), .A(N11799));
MXI2X2 inst_cellmath__25_0_I13777 (.Y(inst_cellmath__25[15]), .A(inst_cellmath__24[14]), .B(inst_cellmath__24[15]), .S0(inst_cellmath__24[47]));
CLKINVX4 inst_cellmath__25_0_I5129 (.Y(N11800), .A(N11799));
NOR2BX1 inst_cellmath__25_0_I2222 (.Y(inst_cellmath__25[0]), .AN(N11807), .B(inst_cellmath__24[0]));
MXI2X1 inst_cellmath__25_0_I2223 (.Y(inst_cellmath__25[1]), .A(inst_cellmath__24[0]), .B(inst_cellmath__24[1]), .S0(N11807));
MX2XL inst_cellmath__25_0_I2224 (.Y(inst_cellmath__25[2]), .A(inst_cellmath__24[1]), .B(inst_cellmath__24[2]), .S0(inst_cellmath__24[47]));
MXI2X1 inst_cellmath__25_0_I2225 (.Y(inst_cellmath__25[3]), .A(inst_cellmath__24[2]), .B(inst_cellmath__24[3]), .S0(N11807));
MXI2X1 inst_cellmath__25_0_I2226 (.Y(inst_cellmath__25[4]), .A(inst_cellmath__24[3]), .B(inst_cellmath__24[4]), .S0(N11807));
MXI2XL inst_cellmath__25_0_I2228 (.Y(inst_cellmath__25[5]), .A(inst_cellmath__24[4]), .B(inst_cellmath__24[5]), .S0(N11800));
MXI2XL inst_cellmath__25_0_I2229 (.Y(inst_cellmath__25[6]), .A(inst_cellmath__24[5]), .B(inst_cellmath__24[6]), .S0(N11800));
MXI2XL inst_cellmath__25_0_I2230 (.Y(inst_cellmath__25[7]), .A(inst_cellmath__24[6]), .B(inst_cellmath__24[7]), .S0(N11800));
MXI2X1 inst_cellmath__25_0_I2231 (.Y(inst_cellmath__25[8]), .A(inst_cellmath__24[7]), .B(inst_cellmath__24[8]), .S0(N11800));
MXI2X1 inst_cellmath__25_0_I2232 (.Y(inst_cellmath__25[9]), .A(inst_cellmath__24[8]), .B(inst_cellmath__24[9]), .S0(N11800));
MXI2X1 inst_cellmath__25_0_I2233 (.Y(inst_cellmath__25[10]), .A(inst_cellmath__24[9]), .B(inst_cellmath__24[10]), .S0(N11800));
MXI2XL inst_cellmath__25_0_I2235 (.Y(inst_cellmath__25[11]), .A(inst_cellmath__24[10]), .B(inst_cellmath__24[11]), .S0(N11801));
MXI2X1 inst_cellmath__25_0_I2236 (.Y(inst_cellmath__25[12]), .A(inst_cellmath__24[11]), .B(inst_cellmath__24[12]), .S0(N11801));
MXI2X1 inst_cellmath__25_0_I2237 (.Y(inst_cellmath__25[13]), .A(inst_cellmath__24[12]), .B(inst_cellmath__24[13]), .S0(N11801));
MXI2X1 inst_cellmath__25_0_I2238 (.Y(inst_cellmath__25[14]), .A(inst_cellmath__24[13]), .B(inst_cellmath__24[14]), .S0(N11801));
MXI2X1 inst_cellmath__25_0_I2240 (.Y(inst_cellmath__25[16]), .A(inst_cellmath__24[15]), .B(inst_cellmath__24[16]), .S0(N11801));
MXI2XL inst_cellmath__25_0_I2242 (.Y(inst_cellmath__25[17]), .A(inst_cellmath__24[16]), .B(inst_cellmath__24[17]), .S0(N11802));
MXI2XL inst_cellmath__25_0_I2243 (.Y(inst_cellmath__25[18]), .A(inst_cellmath__24[17]), .B(inst_cellmath__24[18]), .S0(N11802));
MXI2XL inst_cellmath__25_0_I2244 (.Y(inst_cellmath__25[19]), .A(inst_cellmath__24[18]), .B(inst_cellmath__24[19]), .S0(N11802));
MXI2X1 inst_cellmath__25_0_I2245 (.Y(inst_cellmath__25[20]), .A(inst_cellmath__24[19]), .B(inst_cellmath__24[20]), .S0(N11802));
MXI2X1 inst_cellmath__25_0_I2246 (.Y(inst_cellmath__25[21]), .A(inst_cellmath__24[20]), .B(inst_cellmath__24[21]), .S0(N11802));
XOR2XL cynw_cm_float_mul_ieee_I13779 (.Y(inst_cellmath__24[22]), .A(N3871), .B(N4392));
MXI2X1 inst_cellmath__25_0_I2247 (.Y(inst_cellmath__25[22]), .A(inst_cellmath__24[21]), .B(inst_cellmath__24[22]), .S0(N11802));
MX2XL cynw_cm_float_mul_ieee_I13780 (.Y(inst_cellmath__24[23]), .A(N5096), .B(N3482), .S0(N4392));
INVXL cynw_cm_float_mul_ieee_I13797 (.Y(N11805), .A(N11799));
MXI2X4 inst_cellmath__25_0_I2250 (.Y(inst_cellmath__25[24]), .A(inst_cellmath__24[23]), .B(inst_cellmath__24[24]), .S0(N11805));
MXI2XL inst_cellmath__25_0_I2251 (.Y(inst_cellmath__25[25]), .A(inst_cellmath__24[24]), .B(inst_cellmath__24[25]), .S0(N11805));
MXI2XL inst_cellmath__25_0_I2252 (.Y(inst_cellmath__25[26]), .A(inst_cellmath__24[25]), .B(inst_cellmath__24[26]), .S0(N11805));
MXI2XL inst_cellmath__25_0_I2253 (.Y(inst_cellmath__25[27]), .A(inst_cellmath__24[26]), .B(inst_cellmath__24[27]), .S0(N11805));
MXI2XL inst_cellmath__25_0_I2254 (.Y(inst_cellmath__25[28]), .A(inst_cellmath__24[27]), .B(inst_cellmath__24[28]), .S0(N11805));
MXI2XL inst_cellmath__25_0_I2256 (.Y(inst_cellmath__25[29]), .A(inst_cellmath__24[28]), .B(inst_cellmath__24[29]), .S0(N11803));
MXI2XL inst_cellmath__25_0_I2257 (.Y(inst_cellmath__25[30]), .A(inst_cellmath__24[29]), .B(inst_cellmath__24[30]), .S0(N11803));
MXI2XL inst_cellmath__25_0_I2258 (.Y(inst_cellmath__25[31]), .A(inst_cellmath__24[30]), .B(inst_cellmath__24[31]), .S0(N11803));
MXI2XL inst_cellmath__25_0_I2259 (.Y(inst_cellmath__25[32]), .A(inst_cellmath__24[31]), .B(inst_cellmath__24[32]), .S0(N11803));
MXI2XL inst_cellmath__25_0_I2260 (.Y(inst_cellmath__25[33]), .A(inst_cellmath__24[32]), .B(inst_cellmath__24[33]), .S0(N11803));
MXI2XL inst_cellmath__25_0_I2261 (.Y(inst_cellmath__25[34]), .A(inst_cellmath__24[33]), .B(inst_cellmath__24[34]), .S0(N11803));
MXI2XL inst_cellmath__25_0_I2262 (.Y(inst_cellmath__25[35]), .A(inst_cellmath__24[34]), .B(inst_cellmath__24[35]), .S0(N11804));
MXI2XL inst_cellmath__25_0_I2263 (.Y(inst_cellmath__25[36]), .A(inst_cellmath__24[35]), .B(inst_cellmath__24[36]), .S0(N11804));
MXI2XL inst_cellmath__25_0_I2264 (.Y(inst_cellmath__25[37]), .A(inst_cellmath__24[36]), .B(inst_cellmath__24[37]), .S0(N11804));
MXI2XL inst_cellmath__25_0_I2265 (.Y(inst_cellmath__25[38]), .A(inst_cellmath__24[37]), .B(inst_cellmath__24[38]), .S0(N11804));
MXI2XL inst_cellmath__25_0_I2266 (.Y(inst_cellmath__25[39]), .A(inst_cellmath__24[38]), .B(inst_cellmath__24[39]), .S0(N11804));
MXI2XL inst_cellmath__25_0_I2267 (.Y(inst_cellmath__25[40]), .A(inst_cellmath__24[39]), .B(inst_cellmath__24[40]), .S0(N11804));
MXI2XL inst_cellmath__25_0_I2268 (.Y(inst_cellmath__25[41]), .A(inst_cellmath__24[40]), .B(inst_cellmath__24[41]), .S0(N11806));
MXI2XL inst_cellmath__25_0_I2269 (.Y(inst_cellmath__25[42]), .A(inst_cellmath__24[41]), .B(inst_cellmath__24[42]), .S0(N11806));
MXI2X1 inst_cellmath__25_0_I2270 (.Y(inst_cellmath__25[43]), .A(inst_cellmath__24[42]), .B(inst_cellmath__24[43]), .S0(N11806));
MXI2XL inst_cellmath__25_0_I2273 (.Y(inst_cellmath__25[46]), .A(inst_cellmath__24[45]), .B(inst_cellmath__24[46]), .S0(N11806));
NAND2BXL inst_cellmath__25_0_I2274 (.Y(inst_cellmath__25[47]), .AN(N11807), .B(inst_cellmath__24[46]));
CLKAND2X2 inst_cellmath__45_0_I2275 (.Y(N7548), .A(inst_cellmath__25[25]), .B(inst_cellmath__25[24]));
AND2XL inst_cellmath__45_0_I2276 (.Y(N7516), .A(inst_cellmath__25[26]), .B(inst_cellmath__25[25]));
AND2XL inst_cellmath__45_0_I2277 (.Y(N7440), .A(inst_cellmath__25[27]), .B(inst_cellmath__25[26]));
AND2XL inst_cellmath__45_0_I2278 (.Y(N7497), .A(inst_cellmath__25[28]), .B(inst_cellmath__25[27]));
AND2XL inst_cellmath__45_0_I2279 (.Y(N7424), .A(inst_cellmath__25[29]), .B(inst_cellmath__25[28]));
AND2XL inst_cellmath__45_0_I2280 (.Y(N7478), .A(inst_cellmath__25[30]), .B(inst_cellmath__25[29]));
AND2XL inst_cellmath__45_0_I2281 (.Y(N7538), .A(inst_cellmath__25[31]), .B(inst_cellmath__25[30]));
AND2XL inst_cellmath__45_0_I2282 (.Y(N7463), .A(inst_cellmath__25[31]), .B(inst_cellmath__25[32]));
CLKAND2X2 inst_cellmath__45_0_I2283 (.Y(N7521), .A(inst_cellmath__25[33]), .B(inst_cellmath__25[32]));
AND2XL inst_cellmath__45_0_I2284 (.Y(N7447), .A(inst_cellmath__25[34]), .B(inst_cellmath__25[33]));
CLKAND2X2 inst_cellmath__45_0_I2285 (.Y(N7504), .A(inst_cellmath__25[34]), .B(inst_cellmath__25[35]));
AND2XL inst_cellmath__45_0_I2286 (.Y(N7430), .A(inst_cellmath__25[36]), .B(inst_cellmath__25[35]));
AND2XL inst_cellmath__45_0_I2287 (.Y(N7486), .A(inst_cellmath__25[37]), .B(inst_cellmath__25[36]));
AND2XL inst_cellmath__45_0_I2288 (.Y(N7545), .A(inst_cellmath__25[38]), .B(inst_cellmath__25[37]));
CLKAND2X2 inst_cellmath__45_0_I2289 (.Y(N7469), .A(inst_cellmath__25[39]), .B(inst_cellmath__25[38]));
AND2XL inst_cellmath__45_0_I2290 (.Y(N7527), .A(inst_cellmath__25[40]), .B(inst_cellmath__25[39]));
AND2XL inst_cellmath__45_0_I2291 (.Y(N7452), .A(inst_cellmath__25[41]), .B(inst_cellmath__25[40]));
AND2XL inst_cellmath__45_0_I2292 (.Y(N7513), .A(inst_cellmath__25[42]), .B(inst_cellmath__25[41]));
AND2XL inst_cellmath__45_0_I2293 (.Y(N7435), .A(inst_cellmath__25[43]), .B(inst_cellmath__25[42]));
AND2XL inst_cellmath__45_0_I2294 (.Y(N7493), .A(inst_cellmath__25[43]), .B(inst_cellmath__25[44]));
INVXL inst_cellmath__45_0_I2297 (.Y(inst_cellmath__45[0]), .A(inst_cellmath__25[24]));
NAND2XL inst_cellmath__45_0_I2298 (.Y(N7530), .A(N7516), .B(inst_cellmath__25[24]));
CLKAND2X3 inst_cellmath__45_0_I2299 (.Y(N7500), .A(N7440), .B(N7548));
NAND2XL inst_cellmath__45_0_I2300 (.Y(N7467), .A(N7497), .B(N7516));
AND2XL inst_cellmath__45_0_I2301 (.Y(N7526), .A(N7424), .B(N7440));
NAND2XL inst_cellmath__45_0_I2302 (.Y(N7450), .A(N7478), .B(N7497));
CLKAND2X2 inst_cellmath__45_0_I2303 (.Y(N7511), .A(N7538), .B(N7424));
NAND2XL inst_cellmath__45_0_I2304 (.Y(N7433), .A(N7463), .B(N7478));
AND2XL inst_cellmath__45_0_I2305 (.Y(N7490), .A(N7521), .B(N7538));
NAND2XL inst_cellmath__45_0_I2306 (.Y(N7550), .A(N7447), .B(N7463));
CLKAND2X2 inst_cellmath__45_0_I2307 (.Y(N7473), .A(N7504), .B(N7521));
NAND2XL inst_cellmath__45_0_I2308 (.Y(N7532), .A(N7430), .B(N7447));
AND2XL inst_cellmath__45_0_I2309 (.Y(N7455), .A(N7486), .B(N7504));
NAND2XL inst_cellmath__45_0_I2310 (.Y(N7517), .A(N7545), .B(N7430));
CLKAND2X2 inst_cellmath__45_0_I2311 (.Y(N7441), .A(N7469), .B(N7486));
NAND2XL inst_cellmath__45_0_I2312 (.Y(N7499), .A(N7527), .B(N7545));
AND2XL inst_cellmath__45_0_I2313 (.Y(N7425), .A(N7452), .B(N7469));
NAND2XL inst_cellmath__45_0_I2314 (.Y(N7479), .A(N7513), .B(N7527));
CLKAND2X2 inst_cellmath__45_0_I2315 (.Y(N7540), .A(N7435), .B(N7452));
AND2XL inst_cellmath__45_0_I2316 (.Y(N7522), .A(N7419), .B(N7435));
AND3XL inst_cellmath__45_0_I5366 (.Y(N7506), .A(inst_cellmath__25[47]), .B(inst_cellmath__25[46]), .C(N7419));
INVXL inst_cellmath__45_0_I2318 (.Y(N7546), .A(inst_cellmath__45[0]));
INVXL inst_cellmath__45_0_I2319 (.Y(N7443), .A(N7548));
INVXL inst_cellmath__45_0_I2320 (.Y(N7470), .A(N7530));
NOR2XL inst_cellmath__45_0_I2321 (.Y(N7482), .A(N7467), .B(inst_cellmath__45[0]));
NAND2XL inst_cellmath__45_0_I2322 (.Y(N7437), .A(N7526), .B(N7548));
NOR2XL inst_cellmath__45_0_I2323 (.Y(N7524), .A(N7450), .B(N7530));
NAND2X4 inst_cellmath__45_0_I2324 (.Y(N7495), .A(N7511), .B(N7500));
NOR2XL inst_cellmath__45_0_I2325 (.Y(N7461), .A(N7433), .B(N7467));
NAND2XL inst_cellmath__45_0_I2326 (.Y(N7520), .A(N7490), .B(N7526));
NOR2XL inst_cellmath__45_0_I2327 (.Y(N7446), .A(N7550), .B(N7450));
AND2XL inst_cellmath__45_0_I2328 (.Y(N7503), .A(N7473), .B(N7511));
NOR2XL inst_cellmath__45_0_I2329 (.Y(N7428), .A(N7532), .B(N7433));
NAND2XL inst_cellmath__45_0_I2330 (.Y(N7485), .A(N7455), .B(N7490));
NOR2XL inst_cellmath__45_0_I2331 (.Y(N7543), .A(N7517), .B(N7550));
NAND2X2 inst_cellmath__45_0_I2332 (.Y(N7468), .A(N7473), .B(N7441));
NAND2X1 inst_cellmath__45_0_I2336 (.Y(N7534), .A(N7506), .B(N7540));
INVXL inst_cellmath__45_0_I2337 (.Y(N7481), .A(N7443));
INVXL inst_cellmath__45_0_I2338 (.Y(N7436), .A(N7500));
INVXL inst_cellmath__45_0_I2339 (.Y(N7464), .A(N7482));
INVXL inst_cellmath__45_0_I2340 (.Y(N7494), .A(N7437));
NAND2XL inst_cellmath__45_0_I2342 (.Y(N7475), .A(N7461), .B(N7546));
NOR2XL inst_cellmath__45_0_I2343 (.Y(N7439), .A(N7468), .B(N7495));
NAND4BXL inst_cellmath__45_0_I2344 (.Y(N7505), .AN(N7499), .B(N7493), .C(N7428), .D(N7513));
NAND2XL inst_cellmath__45_0_I2345 (.Y(N7476), .A(N7446), .B(N7470));
NAND2XL inst_cellmath__45_0_I2346 (.Y(N7508), .A(N7503), .B(N7500));
NAND2XL inst_cellmath__45_0_I2347 (.Y(N7537), .A(N7428), .B(N7482));
OR2XL inst_cellmath__45_0_I2348 (.Y(N7432), .A(N7485), .B(N7437));
NAND2XL inst_cellmath__45_0_I2349 (.Y(N7459), .A(N7543), .B(N7524));
NAND4BBXL inst_cellmath__45_0_I2350 (.Y(N7422), .AN(N7499), .BN(N7532), .C(N7546), .D(N7461));
NAND4BXL inst_cellmath__45_0_I2351 (.Y(N7512), .AN(N7520), .B(N7425), .C(N7481), .D(N7455));
NAND4BBXL inst_cellmath__45_0_I2352 (.Y(N7462), .AN(N7479), .BN(N7517), .C(N7470), .D(N7446));
NAND3XL inst_cellmath__45_0_I5250 (.Y(N7484), .A(N7540), .B(N7441), .C(N7503));
NOR2XL inst_cellmath__45_0_I2354 (.Y(N7551), .A(N7436), .B(N7484));
NAND4BXL inst_cellmath__45_0_I2355 (.Y(N7456), .AN(N7485), .B(N7522), .C(N7494), .D(N7425));
NOR3X2 inst_cellmath__45_0_I2358 (.Y(inst_cellmath__45[24]), .A(N7534), .B(N7468), .C(N7495));
XNOR2X1 inst_cellmath__45_0_I2362 (.Y(inst_cellmath__45[4]), .A(N7436), .B(inst_cellmath__25[28]));
XNOR2X1 inst_cellmath__45_0_I2363 (.Y(inst_cellmath__45[5]), .A(N7464), .B(inst_cellmath__25[29]));
XNOR2X1 inst_cellmath__45_0_I2366 (.Y(inst_cellmath__45[8]), .A(N7495), .B(inst_cellmath__25[32]));
XNOR2X1 inst_cellmath__45_0_I2367 (.Y(inst_cellmath__45[9]), .A(N7475), .B(inst_cellmath__25[33]));
NOR2XL inst_cellmath__45_0_I2368 (.Y(N7491), .A(N7520), .B(N7443));
XNOR2X1 inst_cellmath__45_0_I2370 (.Y(inst_cellmath__45[11]), .A(N7476), .B(inst_cellmath__25[35]));
XNOR2X1 inst_cellmath__45_0_I2371 (.Y(inst_cellmath__45[12]), .A(N7508), .B(inst_cellmath__25[36]));
XNOR2X1 inst_cellmath__45_0_I2372 (.Y(inst_cellmath__45[13]), .A(N7537), .B(inst_cellmath__25[37]));
XNOR2X1 inst_cellmath__45_0_I2373 (.Y(inst_cellmath__45[14]), .A(N7432), .B(inst_cellmath__25[38]));
XNOR2X1 inst_cellmath__45_0_I2374 (.Y(inst_cellmath__45[15]), .A(N7459), .B(inst_cellmath__25[39]));
XNOR2X1 inst_cellmath__45_0_I2376 (.Y(inst_cellmath__45[17]), .A(inst_cellmath__25[41]), .B(N7422));
XNOR2X1 inst_cellmath__45_0_I2377 (.Y(inst_cellmath__45[18]), .A(N7512), .B(inst_cellmath__25[42]));
XNOR2X1 inst_cellmath__45_0_I2378 (.Y(inst_cellmath__45[19]), .A(inst_cellmath__25[43]), .B(N7462));
NOR2XL inst_cellmath__45_0_I2380 (.Y(N7429), .A(N7505), .B(N7464));
XNOR2X1 inst_cellmath__45_0_I2382 (.Y(inst_cellmath__45[22]), .A(N7456), .B(inst_cellmath__25[46]));
INVXL inst_cellmath__5_1_I2384 (.Y(N7663), .A(rm[1]));
INVXL inst_cellmath__5_1_I2385 (.Y(N7666), .A(rm[2]));
AND3XL inst_cellmath__5_1_I5252 (.Y(inst_cellmath__5), .A(rm[0]), .B(N7666), .C(N7663));
INVXL inst_cellmath__6_0_I2390 (.Y(N7679), .A(rm[0]));
NAND3XL inst_cellmath__6_0_I2392 (.Y(N7684), .A(rm[1]), .B(N7666), .C(N7679));
NOR2X1 inst_cellmath__34_0_I2404 (.Y(N7749), .A(inst_cellmath__25[0]), .B(inst_cellmath__25[1]));
NOR2X1 inst_cellmath__34_0_I2405 (.Y(N7759), .A(inst_cellmath__25[22]), .B(inst_cellmath__25[21]));
NOR2X1 inst_cellmath__34_0_I2406 (.Y(N7721), .A(inst_cellmath__25[20]), .B(inst_cellmath__25[19]));
NOR2X1 inst_cellmath__34_0_I2407 (.Y(N7731), .A(inst_cellmath__25[18]), .B(inst_cellmath__25[17]));
NOR2X1 inst_cellmath__34_0_I2408 (.Y(N7742), .A(inst_cellmath__25[15]), .B(inst_cellmath__25[16]));
NOR2X1 inst_cellmath__34_0_I2409 (.Y(N7753), .A(inst_cellmath__25[14]), .B(inst_cellmath__25[13]));
NOR2X1 inst_cellmath__34_0_I2410 (.Y(N7763), .A(inst_cellmath__25[12]), .B(inst_cellmath__25[11]));
NOR2XL inst_cellmath__34_0_I2411 (.Y(N7725), .A(inst_cellmath__25[10]), .B(inst_cellmath__25[9]));
NOR2XL inst_cellmath__34_0_I2412 (.Y(N7735), .A(inst_cellmath__25[8]), .B(inst_cellmath__25[7]));
NOR2XL inst_cellmath__34_0_I2413 (.Y(N7746), .A(inst_cellmath__25[6]), .B(inst_cellmath__25[5]));
NOR2XL inst_cellmath__34_0_I2414 (.Y(N7757), .A(inst_cellmath__25[3]), .B(inst_cellmath__25[4]));
NAND2X1 inst_cellmath__34_0_I2416 (.Y(N7729), .A(inst_cellmath__25[2]), .B(N7749));
NAND2X1 inst_cellmath__34_0_I2417 (.Y(N7740), .A(N7759), .B(N7721));
NAND2X2 inst_cellmath__34_0_I2418 (.Y(N7751), .A(N7731), .B(N7742));
NAND2X2 inst_cellmath__34_0_I2419 (.Y(N7761), .A(N7753), .B(N7763));
NAND2XL inst_cellmath__34_0_I2420 (.Y(N7723), .A(N7725), .B(N7735));
NAND2XL inst_cellmath__34_0_I2421 (.Y(N7733), .A(N7757), .B(N7746));
NOR2X1 inst_cellmath__34_0_I2422 (.Y(N7744), .A(N7729), .B(N7740));
NOR2XL inst_cellmath__34_0_I2425 (.Y(N7738), .A(N7723), .B(N7733));
NAND2X1 cynw_cm_float_mul_ieee_I13781 (.Y(N22634), .A(N11788), .B(inst_cellmath__5));
OR2XL cynw_cm_float_mul_ieee_I13782 (.Y(N22643), .A(N11788), .B(N7684));
NAND3XL cynw_cm_float_mul_ieee_I13783 (.Y(N22613), .A(rm[2]), .B(N7663), .C(N7679));
NAND3XL cynw_cm_float_mul_ieee_I13784 (.Y(N22622), .A(N7679), .B(N7663), .C(N7666));
NOR2X6 cynw_cm_float_mul_ieee_I13785 (.Y(N22628), .A(N7751), .B(N7761));
CLKAND2X2 cynw_cm_float_mul_ieee_I13786 (.Y(N22638), .A(N7744), .B(N7738));
NAND2X4 cynw_cm_float_mul_ieee_I13787 (.Y(N22646), .A(N22628), .B(N22638));
NOR2X4 cynw_cm_float_mul_ieee_I13788 (.Y(N22619), .A(inst_cellmath__25[24]), .B(N22646));
NOR2X4 cynw_cm_float_mul_ieee_I13789 (.Y(N22615), .A(N22622), .B(N22619));
NAND2X4 cynw_cm_float_mul_ieee_I13790 (.Y(N22631), .A(N22643), .B(N22634));
BUFX2 cynw_cm_float_mul_ieee_I13791 (.Y(N22617), .A(N22646));
NAND2X4 cynw_cm_float_mul_ieee_I13792 (.Y(N22641), .A(N22617), .B(N22631));
NAND3X8 cynw_cm_float_mul_ieee_I13793 (.Y(N22637), .A(N22613), .B(N22643), .C(N22634));
NOR2X6 cynw_cm_float_mul_ieee_I13794 (.Y(N22614), .A(N22637), .B(N22615));
MX2XL cynw_cm_float_mul_ieee_I14028 (.Y(N22612), .A(inst_cellmath__24[22]), .B(inst_cellmath__24[23]), .S0(N11805));
OAI21X4 cynw_cm_float_mul_ieee_I13799 (.Y(inst_cellmath__44), .A0(N22612), .A1(N22614), .B0(N22641));
INVXL inst_cellmath__30_0_I2448 (.Y(N7857), .A(a_exp[7]));
NOR2XL inst_cellmath__30_0_I2449 (.Y(N7900), .A(a_exp[1]), .B(b_exp[1]));
NAND2XL inst_cellmath__30_0_I2450 (.Y(N7916), .A(a_exp[1]), .B(b_exp[1]));
NOR2XL inst_cellmath__30_0_I2451 (.Y(N7854), .A(a_exp[2]), .B(b_exp[2]));
NAND2XL inst_cellmath__30_0_I2452 (.Y(N7870), .A(a_exp[2]), .B(b_exp[2]));
NOR2XL inst_cellmath__30_0_I2453 (.Y(N7892), .A(a_exp[3]), .B(b_exp[3]));
NAND2XL inst_cellmath__30_0_I2454 (.Y(N7908), .A(a_exp[3]), .B(b_exp[3]));
NOR2XL inst_cellmath__30_0_I2455 (.Y(N7920), .A(a_exp[4]), .B(b_exp[4]));
NAND2XL inst_cellmath__30_0_I2456 (.Y(N7861), .A(a_exp[4]), .B(b_exp[4]));
NOR2XL inst_cellmath__30_0_I2457 (.Y(N7881), .A(a_exp[5]), .B(b_exp[5]));
NAND2XL inst_cellmath__30_0_I2458 (.Y(N7897), .A(a_exp[5]), .B(b_exp[5]));
NOR2XL inst_cellmath__30_0_I2459 (.Y(N7913), .A(a_exp[6]), .B(b_exp[6]));
NAND2XL inst_cellmath__30_0_I2460 (.Y(N7852), .A(a_exp[6]), .B(b_exp[6]));
NOR2XL inst_cellmath__30_0_I2461 (.Y(N7867), .A(b_exp[7]), .B(N7857));
NAND2XL inst_cellmath__30_0_I2462 (.Y(N7888), .A(b_exp[7]), .B(N7857));
OR2XL inst_cellmath__30_0_I2465 (.Y(N7879), .A(b_exp[0]), .B(a_exp[0]));
AOI21XL inst_cellmath__30_0_I2467 (.Y(N7885), .A0(N7870), .A1(N7900), .B0(N7854));
NAND2XL inst_cellmath__30_0_I2468 (.Y(N7903), .A(N7870), .B(N7916));
AOI21XL inst_cellmath__30_0_I2469 (.Y(N7873), .A0(N7861), .A1(N7892), .B0(N7920));
NAND2XL inst_cellmath__30_0_I2470 (.Y(N7894), .A(N7861), .B(N7908));
AOI21XL inst_cellmath__30_0_I2471 (.Y(N7863), .A0(N7852), .A1(N7881), .B0(N7913));
NAND2XL inst_cellmath__30_0_I2472 (.Y(N7882), .A(N7852), .B(N7897));
NAND2XL inst_cellmath__30_0_I2473 (.Y(N7869), .A(N7857), .B(N7867));
NAND2XL inst_cellmath__30_0_I2474 (.Y(N7890), .A(N7857), .B(N7888));
OAI21XL inst_cellmath__30_0_I2475 (.Y(N7859), .A0(N7903), .A1(N7879), .B0(N7885));
INVXL inst_cellmath__30_0_I2476 (.Y(N7891), .A(N7873));
INVXL inst_cellmath__30_0_I2477 (.Y(N7907), .A(N7894));
OAI21XL inst_cellmath__30_0_I2478 (.Y(N7849), .A0(N7882), .A1(N7873), .B0(N7863));
NOR2XL inst_cellmath__30_0_I2479 (.Y(N7865), .A(N7882), .B(N7894));
AOI21XL inst_cellmath__30_0_I2482 (.Y(N7911), .A0(N7865), .A1(N7859), .B0(N7849));
NAND2BXL inst_cellmath__30_0_I2483 (.Y(N7878), .AN(N7900), .B(N7916));
NAND2BXL inst_cellmath__30_0_I2484 (.Y(N7848), .AN(N7854), .B(N7870));
NAND2BXL inst_cellmath__30_0_I2485 (.Y(N7902), .AN(N7892), .B(N7908));
NAND2BXL inst_cellmath__30_0_I2486 (.Y(N7871), .AN(N7920), .B(N7861));
NAND2BXL inst_cellmath__30_0_I2488 (.Y(N7898), .AN(N7913), .B(N7852));
NAND2BXL inst_cellmath__30_0_I2489 (.Y(N7868), .AN(N7867), .B(N7888));
XNOR2X1 inst_cellmath__30_0_I2492 (.Y(inst_cellmath__30[1]), .A(N7879), .B(N7878));
XNOR2X1 inst_cellmath__30_0_I2493 (.Y(inst_cellmath__30[3]), .A(N7859), .B(N7902));
XNOR2X1 inst_cellmath__30_0_I2495 (.Y(inst_cellmath__30[7]), .A(N7911), .B(N7868));
XNOR2X1 inst_cellmath__30_0_I2496 (.Y(N7918), .A(N7848), .B(N7916));
XNOR2X1 inst_cellmath__30_0_I2497 (.Y(N7904), .A(N7848), .B(N7900));
MXI2XL inst_cellmath__30_0_I2498 (.Y(inst_cellmath__30[2]), .A(N7918), .B(N7904), .S0(N7879));
XNOR2X1 inst_cellmath__30_0_I2499 (.Y(N7895), .A(N7871), .B(N7908));
XNOR2X1 inst_cellmath__30_0_I2500 (.Y(N7874), .A(N7871), .B(N7892));
XNOR2X1 inst_cellmath__30_0_I2502 (.Y(N7864), .A(N7898), .B(N7897));
XNOR2X1 inst_cellmath__30_0_I2503 (.Y(N7923), .A(N7898), .B(N7881));
AOI21XL inst_cellmath__31_0_I13898 (.Y(N7875), .A0(N7907), .A1(N7859), .B0(N7891));
MXI2XL inst_cellmath__30_0_I2504 (.Y(inst_cellmath__30[6]), .A(N7864), .B(N7923), .S0(N7875));
XNOR2X1 inst_cellmath__30_0_I2505 (.Y(N7915), .A(N7857), .B(N7888));
XNOR2X1 inst_cellmath__30_0_I2506 (.Y(N7899), .A(N7857), .B(N7867));
MX2XL inst_cellmath__30_0_I2507 (.Y(inst_cellmath__30[8]), .A(N7915), .B(N7899), .S0(N7911));
OAI21XL inst_cellmath__30_0_I2508 (.Y(inst_cellmath__30[9]), .A0(N7890), .A1(N7911), .B0(N7869));
INVXL inst_cellmath__31_0_I13900 (.Y(N22852), .A(N7875));
NOR2BX1 inst_cellmath__31_0_I14031 (.Y(N22875), .AN(N7897), .B(N7881));
INVXL inst_cellmath__31_0_I13902 (.Y(N22848), .A(N22875));
MXI2XL inst_cellmath__31_0_I13903 (.Y(N22871), .A(N22848), .B(N22875), .S0(N22852));
XNOR2X1 inst_cellmath__31_0_I13904 (.Y(inst_cellmath__30[5]), .A(N22875), .B(N22852));
MXI2XL inst_cellmath__31_0_I13905 (.Y(inst_cellmath__30[4]), .A(N7874), .B(N7895), .S0(N7859));
INVXL inst_cellmath__31_0_I13814 (.Y(N22684), .A(b_exp[0]));
INVXL inst_cellmath__31_0_I13815 (.Y(N22696), .A(a_exp[0]));
XOR2XL inst_cellmath__31_0_I13816 (.Y(inst_cellmath__31[0]), .A(N22684), .B(N22696));
NOR2BX1 inst_cellmath__31_0_I2510 (.Y(N8014), .AN(inst_cellmath__30[1]), .B(inst_cellmath__31[0]));
NAND2XL inst_cellmath__31_0_I2511 (.Y(N7994), .A(inst_cellmath__30[2]), .B(N8014));
OR2XL inst_cellmath__31_0_I13906 (.Y(N7998), .A(N7994), .B(inst_cellmath__30[3]));
INVXL inst_cellmath__31_0_I13907 (.Y(N22846), .A(inst_cellmath__30[4]));
NOR2XL inst_cellmath__31_0_I13908 (.Y(N22854), .A(N22846), .B(N7998));
XNOR2X1 inst_cellmath__31_0_I13909 (.Y(N22861), .A(N22846), .B(N7998));
MXI2XL inst_cellmath__31_0_I13911 (.Y(N22869), .A(N22875), .B(N22848), .S0(N7875));
MXI2XL inst_cellmath__31_0_I14032 (.Y(N22865), .A(inst_cellmath__30[5]), .B(N22869), .S0(N22854));
AOI21X2 inst_cellmath__31_0_I13914 (.Y(N22681), .A0(inst_cellmath__45[24]), .A1(inst_cellmath__44), .B0(inst_cellmath__24[47]));
INVX4 inst_cellmath__31_0_I13915 (.Y(inst_cellmath__38), .A(N22681));
MXI2XL inst_cellmath__31_0_I13916 (.Y(N22856), .A(N22846), .B(N22861), .S0(inst_cellmath__38));
MXI2XL inst_cellmath__31_0_I13917 (.Y(N22872), .A(N22871), .B(N22865), .S0(inst_cellmath__38));
NAND2XL inst_cellmath__31_0_I13918 (.Y(N8140), .A(N22856), .B(N22872));
MX2XL inst_cellmath__31_0_I13919 (.Y(inst_cellmath__48[4]), .A(N22846), .B(N22861), .S0(inst_cellmath__38));
NAND2XL node_cs_const1_cs_ii_A_I14134 (.Y(N22987), .A(N22854), .B(inst_cellmath__38));
XOR2XL node_cs_const1_cs_ii_A_I14135 (.Y(inst_cellmath__48[5]), .A(inst_cellmath__30[5]), .B(N22987));
OR2XL inst_cellmath__31_0_I13803 (.Y(inst_cellmath__27), .A(inst_cellmath__14), .B(inst_cellmath__21));
INVXL inst_cellmath__31_0_I2521 (.Y(N7993), .A(inst_cellmath__30[8]));
NAND2XL inst_cellmath__31_0_I2520 (.Y(N8011), .A(inst_cellmath__30[7]), .B(inst_cellmath__30[6]));
XNOR2X1 inst_cellmath__31_0_I2530 (.Y(N8015), .A(N7993), .B(N8011));
NAND2XL hyperpropagate_3_1_A_I5421 (.Y(N11840), .A(inst_cellmath__30[5]), .B(inst_cellmath__30[4]));
NOR2XL hyperpropagate_3_1_A_I5422 (.Y(N8001), .A(N7998), .B(N11840));
MX2XL inst_cellmath__31_0_I2531 (.Y(inst_cellmath__31[8]), .A(N7993), .B(N8015), .S0(N8001));
MX2XL inst_cellmath__48_0_I5158 (.Y(inst_cellmath__48[8]), .A(N7993), .B(inst_cellmath__31[8]), .S0(inst_cellmath__38));
NAND2X1 inst_cellmath__50__50__I2581 (.Y(N8176), .A(inst_cellmath__48[4]), .B(inst_cellmath__48[8]));
INVXL inst_cellmath__31_0_I2523 (.Y(N7991), .A(inst_cellmath__30[7]));
INVXL inst_cellmath__31_0_I2519 (.Y(N8004), .A(inst_cellmath__30[6]));
XNOR2X1 inst_cellmath__31_0_I2528 (.Y(N8018), .A(N7991), .B(N8004));
MX2XL inst_cellmath__31_0_I2529 (.Y(inst_cellmath__31[7]), .A(N7991), .B(N8018), .S0(N8001));
MXI2XL inst_cellmath__48_0_I5040 (.Y(inst_cellmath__48[7]), .A(N7991), .B(inst_cellmath__31[7]), .S0(inst_cellmath__38));
INVXL cynw_cm_float_mul_ieee_I371 (.Y(N1861), .A(inst_cellmath__48[7]));
NAND2X1 inst_cellmath__50__50__I2582 (.Y(N8181), .A(inst_cellmath__48[5]), .B(N1861));
NOR2XL inst_cellmath__50__50__I2586 (.Y(N8187), .A(N8176), .B(N8181));
INVXL inst_cellmath__48_0_I2547 (.Y(N8047), .A(inst_cellmath__30[3]));
XOR2XL inst_cellmath__31_0_I2524 (.Y(inst_cellmath__31[3]), .A(N7994), .B(inst_cellmath__30[3]));
MX2XL inst_cellmath__48_0_I5078 (.Y(inst_cellmath__48[3]), .A(N8047), .B(inst_cellmath__31[3]), .S0(inst_cellmath__38));
MXI2XL inst_cellmath__31_0_I13819 (.Y(N22677), .A(N22696), .B(a_exp[0]), .S0(N22684));
XNOR2X1 inst_cellmath__31_0_I13820 (.Y(inst_cellmath__48[0]), .A(N22681), .B(N22677));
OR2XL inst_cellmath__50__50__I2584 (.Y(N8178), .A(inst_cellmath__48[3]), .B(inst_cellmath__48[0]));
NOR2XL inst_cellmath__31_0_I2522 (.Y(N7990), .A(N7993), .B(N8011));
NAND2XL inst_cellmath__31_0_I2532 (.Y(N8016), .A(N7990), .B(N8001));
XNOR2X1 inst_cellmath__31_0_I2533 (.Y(inst_cellmath__31[9]), .A(inst_cellmath__30[9]), .B(N8016));
MX2XL inst_cellmath__48_0_I5159 (.Y(inst_cellmath__48[9]), .A(inst_cellmath__30[9]), .B(inst_cellmath__31[9]), .S0(inst_cellmath__38));
XNOR2X1 inst_cellmath__31_0_I2512 (.Y(inst_cellmath__31[1]), .A(inst_cellmath__31[0]), .B(inst_cellmath__30[1]));
MX2XL inst_cellmath__48_0_I5154 (.Y(inst_cellmath__48[1]), .A(inst_cellmath__30[1]), .B(inst_cellmath__31[1]), .S0(inst_cellmath__38));
NOR2XL inst_cellmath__50__50__I2579 (.Y(N8188), .A(inst_cellmath__48[9]), .B(inst_cellmath__48[1]));
XOR2XL inst_cellmath__31_0_I2513 (.Y(inst_cellmath__31[2]), .A(N8014), .B(inst_cellmath__30[2]));
MX2XL cynw_cm_float_mul_ieee_I5041 (.Y(N1054), .A(inst_cellmath__30[2]), .B(inst_cellmath__31[2]), .S0(inst_cellmath__38));
XOR2XL inst_cellmath__31_0_I2527 (.Y(inst_cellmath__31[6]), .A(N8001), .B(N8004));
MXI2X1 inst_cellmath__48_0_I5061 (.Y(inst_cellmath__48[6]), .A(N8004), .B(inst_cellmath__31[6]), .S0(inst_cellmath__38));
NOR2XL inst_cellmath__50__50__I2580 (.Y(N8173), .A(inst_cellmath__48[6]), .B(N1054));
NAND2XL inst_cellmath__50__50__I2583 (.Y(N8190), .A(N8188), .B(N8173));
NOR2XL inst_cellmath__50__50__I2585 (.Y(N8183), .A(N8178), .B(N8190));
OR2XL cynw_cm_float_mul_ieee_I5269 (.Y(inst_cellmath__28), .A(inst_cellmath__20), .B(inst_cellmath__13));
OR3XL inst_cellmath__49_1_I5271 (.Y(N8206), .A(inst_cellmath__28), .B(inst_cellmath__27), .C(inst_cellmath__26));
NOR2XL inst_cellmath__49_1_I5163 (.Y(N8212), .A(N8206), .B(inst_cellmath__48[9]));
OAI2BB1X1 inst_cellmath__31_0_I13804 (.Y(N22693), .A0N(N8187), .A1N(N8183), .B0(N8212));
NAND2X1 inst_cellmath__51__49__I2564 (.Y(N8132), .A(inst_cellmath__48[0]), .B(inst_cellmath__48[1]));
NAND2XL inst_cellmath__51__49__I2565 (.Y(N8136), .A(inst_cellmath__48[7]), .B(inst_cellmath__48[6]));
NOR2X2 inst_cellmath__51__49__I2568 (.Y(N8130), .A(N8136), .B(N8132));
NAND2X1 inst_cellmath__51__49__I2567 (.Y(N8127), .A(N1054), .B(inst_cellmath__48[3]));
NOR2X2 inst_cellmath__51__49__I2569 (.Y(N8134), .A(N8140), .B(N8127));
NAND2X2 inst_cellmath__51__49__I2570 (.Y(N8138), .A(N8130), .B(N8134));
DLY1X1 cynw_cm_float_mul_ieee_I2574 (.Y(N8157), .A(inst_cellmath__48[9]));
AOI21X2 inst_cellmath__31_0_I13805 (.Y(N22706), .A0(inst_cellmath__48[8]), .A1(N8138), .B0(N8157));
NOR2X4 inst_cellmath__31_0_I13806 (.Y(N22685), .A(N22706), .B(N22693));
INVX12 inst_cellmath__31_0_I13807 (.Y(inst_cellmath__49), .A(N22685));
NOR2XL cynw_cm_float_mul_ieee_I2597 (.Y(N8228), .A(inst_cellmath__30[8]), .B(inst_cellmath__30[7]));
OR2XL cynw_cm_float_mul_ieee_I2600 (.Y(inst_cellmath__32), .A(inst_cellmath__30[9]), .B(N8228));
OR2XL inst_cellmath__31_0_I13810 (.Y(N469), .A(inst_cellmath__28), .B(inst_cellmath__32));
AND3XL cynw_cm_float_mul_ieee_I5274 (.Y(inst_cellmath__7), .A(rm[0]), .B(rm[1]), .C(N7666));
MXI2XL cynw_cm_float_mul_ieee_I2606 (.Y(N8254), .A(N11788), .B(inst_cellmath__7), .S0(N7684));
MX2XL inst_cellmath__31_0_I13811 (.Y(inst_cellmath__42), .A(N8254), .B(N11788), .S0(inst_cellmath__5));
NOR2BX1 inst_cellmath__31_0_I13812 (.Y(N22689), .AN(inst_cellmath__42), .B(N469));
NOR3XL inst_cellmath__31_0_I13813 (.Y(N22678), .A(N22689), .B(inst_cellmath__27), .C(inst_cellmath__26));
MXI2XL inst_cellmath__31_0_I13817 (.Y(N22682), .A(N22681), .B(inst_cellmath__38), .S0(inst_cellmath__31[0]));
MXI2XL inst_cellmath__31_0_I13818 (.Y(x[23]), .A(N22682), .B(N22678), .S0(inst_cellmath__49));
NOR3BXL inst_cellmath__52_0_I14055 (.Y(N8288), .AN(N469), .B(inst_cellmath__27), .C(inst_cellmath__26));
INVXL inst_cellmath__52_0_I2612 (.Y(N8279), .A(inst_cellmath__48[1]));
INVXL inst_cellmath__52_0_I2613 (.Y(N8285), .A(N1054));
INVXL inst_cellmath__52_0_I2614 (.Y(N8263), .A(inst_cellmath__48[3]));
INVXL inst_cellmath__52_0_I2617 (.Y(N8282), .A(inst_cellmath__48[6]));
MXI2XL inst_cellmath__52_0_I2620 (.Y(x[24]), .A(N8279), .B(N8288), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__52_0_I2621 (.Y(x[25]), .A(N8285), .B(N8288), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__52_0_I2622 (.Y(x[26]), .A(N8263), .B(N8288), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__52_0_I5022 (.Y(x[27]), .A(inst_cellmath__48[4]), .B(N8288), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__52_0_I5023 (.Y(x[28]), .A(inst_cellmath__48[5]), .B(N8288), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__52_0_I2625 (.Y(x[29]), .A(N8282), .B(N8288), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__52_0_I5047 (.Y(x[30]), .A(N1861), .B(N8288), .S0(inst_cellmath__49));
OR4X1 inst_cellmath__47_0_I5275 (.Y(N8319), .A(inst_cellmath__28), .B(inst_cellmath__42), .C(inst_cellmath__26), .D(inst_cellmath__27));
NOR2XL inst_cellmath__47_0_I2629 (.Y(inst_cellmath__47), .A(N8319), .B(inst_cellmath__32));
NOR2XL inst_cellmath__53_U_I2630 (.Y(N8329), .A(inst_cellmath__47), .B(inst_cellmath__26));
MXI2XL inst_cellmath__53_U_I2631 (.Y(N8324), .A(inst_cellmath__25[46]), .B(inst_cellmath__45[22]), .S0(inst_cellmath__44));
MXI2XL inst_cellmath__53_U_I2632 (.Y(x[22]), .A(N8324), .B(N8329), .S0(inst_cellmath__49));
AND2XL inst_cellmath__53_M_I2635 (.Y(N8472), .A(b_man[0]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2636 (.Y(N8348), .A(b_man[1]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2637 (.Y(N8447), .A(b_man[2]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2638 (.Y(N8541), .A(b_man[3]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2639 (.Y(N8417), .A(b_man[4]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2640 (.Y(N8512), .A(b_man[5]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2641 (.Y(N8390), .A(b_man[6]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2642 (.Y(N8484), .A(b_man[7]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2643 (.Y(N8361), .A(b_man[8]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2644 (.Y(N8458), .A(b_man[9]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2645 (.Y(N8554), .A(b_man[10]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2646 (.Y(N8430), .A(b_man[11]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2647 (.Y(N8525), .A(b_man[12]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2648 (.Y(N8401), .A(b_man[13]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2649 (.Y(N8495), .A(b_man[14]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2650 (.Y(N8373), .A(b_man[15]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2651 (.Y(N8468), .A(b_man[16]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2652 (.Y(N8342), .A(b_man[17]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2653 (.Y(N8442), .A(b_man[18]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2654 (.Y(N8536), .A(b_man[19]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2655 (.Y(N8411), .A(b_man[20]), .B(inst_cellmath__22));
AND2XL inst_cellmath__53_M_I2656 (.Y(N8507), .A(b_man[21]), .B(inst_cellmath__22));
MX2XL inst_cellmath__53_M_I2659 (.Y(N8384), .A(N8472), .B(a_man[0]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2660 (.Y(N8434), .A(N8348), .B(a_man[1]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2661 (.Y(N8479), .A(N8447), .B(a_man[2]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2662 (.Y(N8529), .A(N8541), .B(a_man[3]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2663 (.Y(N8354), .A(N8417), .B(a_man[4]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2664 (.Y(N8404), .A(N8512), .B(a_man[5]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2665 (.Y(N8454), .A(N8390), .B(a_man[6]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2666 (.Y(N8499), .A(N8484), .B(a_man[7]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2667 (.Y(N8549), .A(N8361), .B(a_man[8]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2668 (.Y(N8377), .A(N8458), .B(a_man[9]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2669 (.Y(N8423), .A(N8554), .B(a_man[10]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2670 (.Y(N8470), .A(N8430), .B(a_man[11]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2671 (.Y(N8519), .A(N8525), .B(a_man[12]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2672 (.Y(N8346), .A(N8401), .B(a_man[13]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2673 (.Y(N8396), .A(N8495), .B(a_man[14]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2674 (.Y(N8446), .A(N8373), .B(a_man[15]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2675 (.Y(N8489), .A(N8468), .B(a_man[16]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2676 (.Y(N8539), .A(N8342), .B(a_man[17]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2677 (.Y(N8368), .A(N8442), .B(a_man[18]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2678 (.Y(N8415), .A(N8536), .B(a_man[19]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2679 (.Y(N8463), .A(N8411), .B(a_man[20]), .S0(inst_cellmath__15));
MX2XL inst_cellmath__53_M_I2680 (.Y(N8511), .A(N8507), .B(a_man[21]), .S0(inst_cellmath__15));
INVXL inst_cellmath__53_M_I2683 (.Y(N8545), .A(inst_cellmath__26));
INVXL inst_cellmath__53_M_I2684 (.Y(N8416), .A(N8545));
MXI2XL inst_cellmath__53_M_I2685 (.Y(N8337), .A(inst_cellmath__47), .B(N8384), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2686 (.Y(N8388), .A(inst_cellmath__47), .B(N8434), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2687 (.Y(N8439), .A(inst_cellmath__47), .B(N8479), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2688 (.Y(N8483), .A(inst_cellmath__47), .B(N8529), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2689 (.Y(N8533), .A(inst_cellmath__47), .B(N8354), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2690 (.Y(N8360), .A(inst_cellmath__47), .B(N8404), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2691 (.Y(N8408), .A(inst_cellmath__47), .B(N8454), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2692 (.Y(N8457), .A(inst_cellmath__47), .B(N8499), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2693 (.Y(N8504), .A(inst_cellmath__47), .B(N8549), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2694 (.Y(N8553), .A(inst_cellmath__47), .B(N8377), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2695 (.Y(N8381), .A(inst_cellmath__47), .B(N8423), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2696 (.Y(N8429), .A(inst_cellmath__47), .B(N8470), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2697 (.Y(N8474), .A(inst_cellmath__47), .B(N8519), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2698 (.Y(N8522), .A(inst_cellmath__47), .B(N8346), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2699 (.Y(N8351), .A(inst_cellmath__47), .B(N8396), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2700 (.Y(N8400), .A(inst_cellmath__47), .B(N8446), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2701 (.Y(N8450), .A(inst_cellmath__47), .B(N8489), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2702 (.Y(N8494), .A(inst_cellmath__47), .B(N8539), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2703 (.Y(N8543), .A(inst_cellmath__47), .B(N8368), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2704 (.Y(N8371), .A(inst_cellmath__47), .B(N8415), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2705 (.Y(N8420), .A(inst_cellmath__47), .B(N8463), .S0(N8416));
MXI2XL inst_cellmath__53_M_I2706 (.Y(N8467), .A(inst_cellmath__47), .B(N8511), .S0(N8416));
INVXL inst_cellmath__53_M_I2707 (.Y(N8524), .A(inst_cellmath__44));
INVXL inst_cellmath__53_M_I2708 (.Y(N8347), .A(N8524));
MXI2XL inst_cellmath__53_M_I2709 (.Y(N8515), .A(inst_cellmath__25[24]), .B(inst_cellmath__45[0]), .S0(N8347));
NAND2XL node_cs_const1_cs_ii_A_I5423 (.Y(N11847), .A(N7546), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5424 (.Y(N8341), .A(inst_cellmath__25[25]), .B(N11847));
NAND2XL node_cs_const1_cs_ii_A_I5425 (.Y(N11854), .A(N7481), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5426 (.Y(N8391), .A(inst_cellmath__25[26]), .B(N11854));
NAND2XL node_cs_const1_cs_ii_A_I5427 (.Y(N11861), .A(N7470), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5428 (.Y(N8440), .A(inst_cellmath__25[27]), .B(N11861));
MXI2XL inst_cellmath__53_M_I2713 (.Y(N8486), .A(inst_cellmath__25[28]), .B(inst_cellmath__45[4]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2714 (.Y(N8535), .A(inst_cellmath__25[29]), .B(inst_cellmath__45[5]), .S0(N8347));
NAND2XL node_cs_const1_cs_ii_A_I5429 (.Y(N11868), .A(N7494), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5430 (.Y(N8363), .A(inst_cellmath__25[30]), .B(N11868));
NAND2XL node_cs_const1_cs_ii_A_I5431 (.Y(N11875), .A(N7524), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5432 (.Y(N8410), .A(inst_cellmath__25[31]), .B(N11875));
MXI2XL inst_cellmath__53_M_I2717 (.Y(N8459), .A(inst_cellmath__25[32]), .B(inst_cellmath__45[8]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2718 (.Y(N8506), .A(inst_cellmath__25[33]), .B(inst_cellmath__45[9]), .S0(N8347));
NAND2XL node_cs_const1_cs_ii_A_I5433 (.Y(N11882), .A(N7491), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5434 (.Y(N8556), .A(inst_cellmath__25[34]), .B(N11882));
MXI2XL inst_cellmath__53_M_I2720 (.Y(N8383), .A(inst_cellmath__25[35]), .B(inst_cellmath__45[11]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2721 (.Y(N8432), .A(inst_cellmath__25[36]), .B(inst_cellmath__45[12]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2722 (.Y(N8477), .A(inst_cellmath__25[37]), .B(inst_cellmath__45[13]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2723 (.Y(N8526), .A(inst_cellmath__25[38]), .B(inst_cellmath__45[14]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2724 (.Y(N8352), .A(inst_cellmath__25[39]), .B(inst_cellmath__45[15]), .S0(N8347));
NAND2XL node_cs_const1_cs_ii_A_I5435 (.Y(N11889), .A(N7439), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5436 (.Y(N8403), .A(inst_cellmath__25[40]), .B(N11889));
MXI2XL inst_cellmath__53_M_I2726 (.Y(N8452), .A(inst_cellmath__25[41]), .B(inst_cellmath__45[17]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2727 (.Y(N8497), .A(inst_cellmath__25[42]), .B(inst_cellmath__45[18]), .S0(N8347));
MXI2XL inst_cellmath__53_M_I2728 (.Y(N8547), .A(inst_cellmath__25[43]), .B(inst_cellmath__45[19]), .S0(N8347));
NAND2XL node_cs_const1_cs_ii_A_I5437 (.Y(N11896), .A(N7551), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5438 (.Y(N8374), .A(inst_cellmath__25[44]), .B(N11896));
NAND2XL node_cs_const1_cs_ii_A_I5439 (.Y(N11903), .A(N7429), .B(N8347));
XOR2XL node_cs_const1_cs_ii_A_I5440 (.Y(N8421), .A(inst_cellmath__25[45]), .B(N11903));
MXI2XL inst_cellmath__53_M_I2733 (.Y(x[0]), .A(N8515), .B(N8337), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2734 (.Y(x[1]), .A(N8341), .B(N8388), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2735 (.Y(x[2]), .A(N8391), .B(N8439), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2736 (.Y(x[3]), .A(N8440), .B(N8483), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2737 (.Y(x[4]), .A(N8486), .B(N8533), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2738 (.Y(x[5]), .A(N8535), .B(N8360), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2739 (.Y(x[6]), .A(N8363), .B(N8408), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2740 (.Y(x[7]), .A(N8410), .B(N8457), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2741 (.Y(x[8]), .A(N8459), .B(N8504), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2742 (.Y(x[9]), .A(N8506), .B(N8553), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2743 (.Y(x[10]), .A(N8556), .B(N8381), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2744 (.Y(x[11]), .A(N8383), .B(N8429), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2745 (.Y(x[12]), .A(N8432), .B(N8474), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2746 (.Y(x[13]), .A(N8477), .B(N8522), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2747 (.Y(x[14]), .A(N8526), .B(N8351), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2748 (.Y(x[15]), .A(N8352), .B(N8400), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2749 (.Y(x[16]), .A(N8403), .B(N8450), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2750 (.Y(x[17]), .A(N8452), .B(N8494), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2751 (.Y(x[18]), .A(N8497), .B(N8543), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2752 (.Y(x[19]), .A(N8547), .B(N8371), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2753 (.Y(x[20]), .A(N8374), .B(N8420), .S0(inst_cellmath__49));
MXI2XL inst_cellmath__53_M_I2754 (.Y(x[21]), .A(N8421), .B(N8467), .S0(inst_cellmath__49));
assign inst_cellmath__24[44] = 1'B0;
assign inst_cellmath__25[23] = 1'B0;
assign inst_cellmath__30[0] = 1'B0;
assign inst_cellmath__31[4] = 1'B0;
assign inst_cellmath__31[5] = 1'B0;
assign inst_cellmath__45[1] = 1'B0;
assign inst_cellmath__45[2] = 1'B0;
assign inst_cellmath__45[3] = 1'B0;
assign inst_cellmath__45[6] = 1'B0;
assign inst_cellmath__45[7] = 1'B0;
assign inst_cellmath__45[10] = 1'B0;
assign inst_cellmath__45[16] = 1'B0;
assign inst_cellmath__45[20] = 1'B0;
assign inst_cellmath__45[21] = 1'B0;
assign inst_cellmath__45[23] = 1'B0;
assign inst_cellmath__48[2] = 1'B0;
endmodule

/* CADENCE  ubD4Sg7Wqhw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



