/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:09 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3784,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3850,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4000,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4017,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4033,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4059,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4784,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4850,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4866,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4921,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5000,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5017,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5059,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22921,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22987;
wire N10691,N10693,N10698,N10700,N10702,N10705,N10707 
	,N10712,N10714,N10719,N10721,N10726,N10728,N10733,N10735 
	,N10740,N10742,N10747,N10749,N10754,N10756,N10761,N10763 
	,N10768,N10770,N10775,N10777,N10782,N10784,N10789,N10791 
	,N10796,N10798,N10803,N10805,N10810,N10812,N10817,N10819 
	,N10824,N10826,N10831,N10833,N10838,N10840,N10847,N10852 
	,N10854,N10861,N10868,N10875,N10882,N10889,N10894,N10896 
	,N10901,N10903,N11175,N11176,N11177,N11178,N11179,N11180 
	,N11181,N11189,N11190,N11217,N11222;
reg x_reg_23__retimed_I6214_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6214_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22682;
	end
assign N10903 = x_reg_23__retimed_I6214_QOUT;
reg x_reg_23__retimed_I6213_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I6213_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22678;
	end
assign N10901 = x_reg_23__retimed_I6213_QOUT;
reg x_reg_22__retimed_I6211_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6211_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8324;
	end
assign N10896 = x_reg_22__retimed_I6211_QOUT;
reg x_reg_22__retimed_I6210_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6210_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8329;
	end
assign N10894 = x_reg_22__retimed_I6210_QOUT;
reg x_reg_24__retimed_I6208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I6208_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8279;
	end
assign N10889 = x_reg_24__retimed_I6208_QOUT;
reg x_reg_25__retimed_I6205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_25__retimed_I6205_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8285;
	end
assign N10882 = x_reg_25__retimed_I6205_QOUT;
reg x_reg_26__retimed_I6202_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__retimed_I6202_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8263;
	end
assign N10875 = x_reg_26__retimed_I6202_QOUT;
reg x_reg_27__retimed_I6199_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__retimed_I6199_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[4];
	end
assign N10868 = x_reg_27__retimed_I6199_QOUT;
reg x_reg_28__retimed_I6196_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__retimed_I6196_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[5];
	end
assign N10861 = x_reg_28__retimed_I6196_QOUT;
reg x_reg_29__retimed_I6193_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__retimed_I6193_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8282;
	end
assign N10854 = x_reg_29__retimed_I6193_QOUT;
reg x_reg_29__retimed_I6192_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__retimed_I6192_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8288;
	end
assign N10852 = x_reg_29__retimed_I6192_QOUT;
reg x_reg_30__retimed_I6190_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__retimed_I6190_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861;
	end
assign N10847 = x_reg_30__retimed_I6190_QOUT;
reg x_reg_0__retimed_I6187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I6187_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8515;
	end
assign N10840 = x_reg_0__retimed_I6187_QOUT;
reg x_reg_0__retimed_I6186_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I6186_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8337;
	end
assign N10838 = x_reg_0__retimed_I6186_QOUT;
reg x_reg_1__retimed_I6184_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I6184_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8341;
	end
assign N10833 = x_reg_1__retimed_I6184_QOUT;
reg x_reg_1__retimed_I6183_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I6183_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8388;
	end
assign N10831 = x_reg_1__retimed_I6183_QOUT;
reg x_reg_2__retimed_I6181_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I6181_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8391;
	end
assign N10826 = x_reg_2__retimed_I6181_QOUT;
reg x_reg_2__retimed_I6180_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I6180_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8439;
	end
assign N10824 = x_reg_2__retimed_I6180_QOUT;
reg x_reg_3__retimed_I6178_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I6178_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8440;
	end
assign N10819 = x_reg_3__retimed_I6178_QOUT;
reg x_reg_3__retimed_I6177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I6177_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8483;
	end
assign N10817 = x_reg_3__retimed_I6177_QOUT;
reg x_reg_4__retimed_I6175_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I6175_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8486;
	end
assign N10812 = x_reg_4__retimed_I6175_QOUT;
reg x_reg_4__retimed_I6174_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I6174_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8533;
	end
assign N10810 = x_reg_4__retimed_I6174_QOUT;
reg x_reg_5__retimed_I6172_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I6172_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8535;
	end
assign N10805 = x_reg_5__retimed_I6172_QOUT;
reg x_reg_5__retimed_I6171_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I6171_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8360;
	end
assign N10803 = x_reg_5__retimed_I6171_QOUT;
reg x_reg_6__retimed_I6169_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I6169_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8363;
	end
assign N10798 = x_reg_6__retimed_I6169_QOUT;
reg x_reg_6__retimed_I6168_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I6168_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8408;
	end
assign N10796 = x_reg_6__retimed_I6168_QOUT;
reg x_reg_7__retimed_I6166_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I6166_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8410;
	end
assign N10791 = x_reg_7__retimed_I6166_QOUT;
reg x_reg_7__retimed_I6165_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I6165_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8457;
	end
assign N10789 = x_reg_7__retimed_I6165_QOUT;
reg x_reg_8__retimed_I6163_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I6163_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8459;
	end
assign N10784 = x_reg_8__retimed_I6163_QOUT;
reg x_reg_8__retimed_I6162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I6162_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8504;
	end
assign N10782 = x_reg_8__retimed_I6162_QOUT;
reg x_reg_9__retimed_I6160_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I6160_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8506;
	end
assign N10777 = x_reg_9__retimed_I6160_QOUT;
reg x_reg_9__retimed_I6159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I6159_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8553;
	end
assign N10775 = x_reg_9__retimed_I6159_QOUT;
reg x_reg_10__retimed_I6157_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I6157_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8556;
	end
assign N10770 = x_reg_10__retimed_I6157_QOUT;
reg x_reg_10__retimed_I6156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I6156_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8381;
	end
assign N10768 = x_reg_10__retimed_I6156_QOUT;
reg x_reg_11__retimed_I6154_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6154_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8383;
	end
assign N10763 = x_reg_11__retimed_I6154_QOUT;
reg x_reg_11__retimed_I6153_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6153_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8429;
	end
assign N10761 = x_reg_11__retimed_I6153_QOUT;
reg x_reg_12__retimed_I6151_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I6151_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8432;
	end
assign N10756 = x_reg_12__retimed_I6151_QOUT;
reg x_reg_12__retimed_I6150_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I6150_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8474;
	end
assign N10754 = x_reg_12__retimed_I6150_QOUT;
reg x_reg_13__retimed_I6148_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I6148_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8477;
	end
assign N10749 = x_reg_13__retimed_I6148_QOUT;
reg x_reg_13__retimed_I6147_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I6147_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8522;
	end
assign N10747 = x_reg_13__retimed_I6147_QOUT;
reg x_reg_14__retimed_I6145_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6145_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8526;
	end
assign N10742 = x_reg_14__retimed_I6145_QOUT;
reg x_reg_14__retimed_I6144_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6144_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8351;
	end
assign N10740 = x_reg_14__retimed_I6144_QOUT;
reg x_reg_15__retimed_I6142_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I6142_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8352;
	end
assign N10735 = x_reg_15__retimed_I6142_QOUT;
reg x_reg_15__retimed_I6141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I6141_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8400;
	end
assign N10733 = x_reg_15__retimed_I6141_QOUT;
reg x_reg_16__retimed_I6139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I6139_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8403;
	end
assign N10728 = x_reg_16__retimed_I6139_QOUT;
reg x_reg_16__retimed_I6138_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I6138_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8450;
	end
assign N10726 = x_reg_16__retimed_I6138_QOUT;
reg x_reg_17__retimed_I6136_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6136_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8452;
	end
assign N10721 = x_reg_17__retimed_I6136_QOUT;
reg x_reg_17__retimed_I6135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6135_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8494;
	end
assign N10719 = x_reg_17__retimed_I6135_QOUT;
reg x_reg_18__retimed_I6133_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I6133_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8497;
	end
assign N10714 = x_reg_18__retimed_I6133_QOUT;
reg x_reg_18__retimed_I6132_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I6132_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8543;
	end
assign N10712 = x_reg_18__retimed_I6132_QOUT;
reg x_reg_19__retimed_I6130_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6130_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8547;
	end
assign N10707 = x_reg_19__retimed_I6130_QOUT;
reg x_reg_19__retimed_I6129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6129_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8371;
	end
assign N10705 = x_reg_19__retimed_I6129_QOUT;
reg x_reg_20__retimed_I6128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6128_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49;
	end
assign N10702 = x_reg_20__retimed_I6128_QOUT;
assign N11190 = !N10702;
assign N11189 = !N10702;
assign N11181 = !N11190;
assign N11180 = !N11189;
assign N11179 = !N11189;
assign N11178 = !N11189;
assign N11177 = !N11189;
assign N11176 = !N11189;
assign N11175 = !N11189;
reg x_reg_20__retimed_I6127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6127_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8374;
	end
assign N10700 = x_reg_20__retimed_I6127_QOUT;
reg x_reg_20__retimed_I6126_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6126_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8420;
	end
assign N10698 = x_reg_20__retimed_I6126_QOUT;
reg x_reg_21__retimed_I6124_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6124_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8421;
	end
assign N10693 = x_reg_21__retimed_I6124_QOUT;
reg x_reg_21__retimed_I6123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6123_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8467;
	end
assign N10691 = x_reg_21__retimed_I6123_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 = !b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4362 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666 = !a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4063 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 = !b_man[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144 = !a_man[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3187 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3557, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3106} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4063} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4362} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3187};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 = !b_man[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672 = !a_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3808 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4090 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133 = !a_man[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4967 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 = !b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4984 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5097, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4643} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4967} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4090} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4984};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3932, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3483} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3808} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3557} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4643};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4977 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4081 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 = !b_man[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4635 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184 = !a_man[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3157 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3464 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3181, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4795} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3157} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4635} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3464};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4461, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4010} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4081} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4977} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3181};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3178 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4351 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4072 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4084, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3635} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4351} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3178} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4072};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3453 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4626 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4340 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4876, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4427} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4626} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3453} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4340};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 = !b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4909 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715 = !a_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4326 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3735 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3976, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3526} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4326} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4909} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3735};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4991, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4538} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3976} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4876} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4795};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3285, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4912} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4084} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3106} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4991};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4461} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3483} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3285};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 = !b_man[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3116 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176 = !a_man[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3425 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4012 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3862, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3412} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3425} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3116} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4012};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3165 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3727 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4901 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4618 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4763, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4313} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4901} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3727} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4618};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3712, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3256} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3165} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3862} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4763};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4332 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3443 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 = !b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3387 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 = !a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4590 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4278 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4920, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4469} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4590} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3387} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4278};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3599, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3147} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4332} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4920};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4611, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4158} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3526} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4427} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3599};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3822, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3364} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3635} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3712} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4611};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4010} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3822} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4912};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4607 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3716 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3433 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4653, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4201} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3716} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4607} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3433};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4001 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3103 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4893 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3755, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3295} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3103} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4001} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4893};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4503, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4054} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3755} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4653} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3412};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4267 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3375 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3094 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3903, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3456} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3375} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4267} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3094};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 = !b_man[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3662 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232 = !a_man[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3689 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4557 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5074, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4620} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3689} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3662} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4557};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4883 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3992 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3707 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4806, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4356} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3992} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4883} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3707};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3493, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5105} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5074} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3903} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4806};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3332, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4952} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3493} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3147};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3446, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5066} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4503} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3256} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3332};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4538} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3446} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3364};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4393, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3940} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4469} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3295} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4201};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3085 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4258 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3983 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4060, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3610} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4258} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3085} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3983};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4547, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4095} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4060} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4620} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3456};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 = !b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3935 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758 = !a_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4854 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4824 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4321, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3872} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4854} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3935} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4824};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4598 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4549 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3651 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3366 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3156, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4772} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3651} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4549} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3366};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3643, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3189} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4598} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4321} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3156};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3225, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4841} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3643} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4547} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5105};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4236, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3790} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4393} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4054} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3225};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4158} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4236} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5066};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3697 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4873 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 = !b_man[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4203 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220 = !a_man[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3951 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5099 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4739, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4289} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3951} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4203} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5099};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4962, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4513} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4873} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3697} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4739};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3356 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4536 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4250 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4480, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4030} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4536} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3356} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4250};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4814 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3926 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3641 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3574, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3122} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3926} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4814} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3641};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3971 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5144 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4864 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3306, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4929} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5144} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3971} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4864};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3800, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3341} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3574} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4480} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3306};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3377, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4998} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4356} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4962} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3800};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4696, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4245} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3872} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4772} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3610};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4280, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3830} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3189} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4696} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4095};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4128, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3678} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3377} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3940} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4280};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4952} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4128} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3790};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5089 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4196 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3915 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3088, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4703} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4196} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5089} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3915};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 = !b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4484 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 = !a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5116 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3298 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4253, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3806} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5116} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4484} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3298};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3634 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4805 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4526 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3994, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3542} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4805} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3634} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4526};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4209, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3764} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4253} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3088} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3994};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4243 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3348 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5135 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4896, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4446} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3348} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4243} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5135};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5112, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4663} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4896} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4289} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3122};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3534, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3081} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4209} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4513} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5112};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 = !b_man[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4751 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273 = !a_man[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4213 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3576 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4939, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4489} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4751} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3576};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3961 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4183 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4476 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3290 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3775, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3316} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4476} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4183} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3290};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3730, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3271} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3961} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4939} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3775};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3950, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3503} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4030} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4929} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3730};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4439, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3986} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3341} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3950} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4245};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3114, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4728} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3534} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4998} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4439};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4841} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3114} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3678};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3467, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5082} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4703} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3542} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4446};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4518 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3626 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3340 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3512, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5121} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3626} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4518} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3340};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3905 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5081 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4797 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4673, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4219} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5081} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3905} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4797};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4628, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4176} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4673} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3512} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3806};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4849, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4403} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4628} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3467} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3764};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5071 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3282 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4175 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4455, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4004} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3282} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5071} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4175};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4741 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3569 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4464 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3550, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3098} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3569} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4741} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4464};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4787 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3893 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3617 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3280, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4904} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3893} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4787} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3617};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3241, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4860} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3550} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4455} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3280};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5125 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4234 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 = !b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5029 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801 = !a_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3307 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3852 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4712, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3307} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5029} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3852};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4410, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3960} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4234} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5125} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4712};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3326 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4508 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4222 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4186, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3740} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4508} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3326} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4222};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4142, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3692} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4186} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4489} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3316};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4366, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3913} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4410} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3241} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4142};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3685, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3234} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4663} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3503} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4366};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3264, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4884} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4849} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3081} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3685};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3830} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3264} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4728};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3843 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5019 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4731 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4499, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4047} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3843} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5019} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4731};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 = !b_man[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3231 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260 = !a_man[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4483 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4125 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3593, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3140} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4483} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3231} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4125};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4453 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3559 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3273 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3324, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4948} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3559} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3273} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4453};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5090, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4637} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3593} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3324};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5049, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4597} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4219} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5121} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5090};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3197, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4816} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3271} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4176} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5049};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3608 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4779 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4501 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5133, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4681} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4779} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3608} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4501};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5065 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4169 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3885 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4229, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3784} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4169} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5065} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3885};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3924, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3476} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4229} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5133} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4262};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4826, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4376} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4904} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4004} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3098};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3881, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3428} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3924} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3960} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4826};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4103, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3653} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5082} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3881} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3913};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4589, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4135} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3197} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4403} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4103};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3986} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4589} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4884};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 = !b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3508 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792 = !a_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3579 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4400 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3638, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3184} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3508} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4400};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3317 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5009 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4114 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3223 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4543, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4086} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4114} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5009} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3223};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3969, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3521} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3317} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4543};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3263 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4160 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4445 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4274, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3825} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4160} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3263} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4445};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4724 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3832 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3549 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3368, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4994} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3832} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4724} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3549};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3876 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5055 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4770 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3110, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4722} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5055} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3876} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4770};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4869, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4420} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3368} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4274} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3110};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3664, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3207} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3740} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3969} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4869};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4780, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4328} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4860} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3692} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3664};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3705, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3250} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3140} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4948} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4047};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4493 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3597 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 = !b_man[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3781 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318 = !a_man[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4740 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4668 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4843, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4397} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4740} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3781} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4668};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4014, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3561} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4493} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4843};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4605, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4153} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3784} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4681} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4014};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4564, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4112} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3705} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4637} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4605};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3621, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3163} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4564} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3428};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5006, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4555} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4780} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4816} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3621};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3234} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5006} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4135};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4760 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3869 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3587 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3150, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4767} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3869} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4760} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3587};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4150 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3254 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5047 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4316, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3867} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3254} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4150} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5047};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3749, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3288} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4316} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3150} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3184};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5001 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4105 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3824 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4581, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4131} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5001} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4105} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3824};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4389 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3501 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3212 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3681, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3228} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3501} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3212} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4389};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4714 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3541 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4436 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3415, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5036} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4436} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3541} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4714};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4915, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4465} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3681} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4581} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3415};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3439, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5059} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4915} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3749} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3521};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3397, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5017} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3476} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4376} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3439};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4646, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4197} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4086} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4994} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3825};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4339, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3889} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4646} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4420} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3250};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4299, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3848} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3207} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4339} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4112};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4520, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4067} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3397} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4328} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4299};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3653} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4520} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4555};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 = !b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4052 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845 = !a_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3842 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4942 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3084, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4699} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3842} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4052} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4942};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4098 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3202 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4378 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4888, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4442} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3202} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4098} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4378};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4660 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3774 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3490 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3990, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3537} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3774} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4660} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3490};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4056, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3602} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4888} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3084} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3990};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3245 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3536 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4426 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4623, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4170} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4426} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3245} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3536};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3814 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4993 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4705 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3726, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3267} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4993} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3814} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4705};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5039 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4141 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3859 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3459, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5078} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4141} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5039} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3859};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4956, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4507} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3726} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4623} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3459};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3488, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5100} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4722} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4056} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4956};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3793, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3337} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4397} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3228} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4131};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4386, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3933} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3561} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3793} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4465};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3174, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4789} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3488} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4153} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4386};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4690, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4239} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4767} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3867} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5036};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3217, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4835} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4690} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3288} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4197};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4077, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3628} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5059} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3889};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3131, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4749} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5017} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4077};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3163} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3131} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4067};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5003, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4551} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4442} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4170} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3267};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4431, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3980} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5003} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3602} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4507};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4982 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3191 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4088 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3125, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4743} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3191} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4982} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4088};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3528 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4695 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3805 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4033, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3578} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4695} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3528} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3805};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4368 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3478 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4650 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4294, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3841} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3478} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4368} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4650};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3193, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4808} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4033} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3125} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4294};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4750 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4043 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4935 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3760 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3392, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5011} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4935} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4043} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3760};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299 = !a_man[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5012 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3146 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737 = !b_man[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11793 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11793;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4320 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4559, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4107} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3146} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5012} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4320};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4361, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3909} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3392} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4750} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4559};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3238 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4417 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4133 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4934, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4482} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4417} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4133} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3238};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4096, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3647} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4699} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4934} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3537};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3529, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5143} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4361} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3193} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4096};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4123, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3673} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3529} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4431} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5100};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3851 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5031 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835 = !a_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4104 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 = !b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4596 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3420 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5124, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4675} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4596} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4104} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3420};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3768, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3309} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5031} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3851} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5124};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4927 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3752 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4640 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4863, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4413} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4927} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3752} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4640};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3138 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4312 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4036 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3963, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3515} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4312} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3138} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4036};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4359 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3183 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3469 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3696, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3244} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3183} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4359} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3469};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4666, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4212} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3963} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4863} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3696};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3833, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3379} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3768} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5078} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4666};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3258, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4878} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4239} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3833} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3337};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5027, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4572} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3258} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3933} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4835};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4983, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4789} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4123} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5027};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3848} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4983} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4749};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4685 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3519 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4409 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3432, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5051} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3519} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4685} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4409};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4079 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4973 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3797 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4600, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4147} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4973} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4079} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3797};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4124 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3230 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5021 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4331, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3884} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3230} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4124} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5021};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3507, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5115} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4600} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3432} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4331};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4729, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4284} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3507} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3909} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4808};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3237, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4853} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4743} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3578} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4482};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4406, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3953} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5011} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4107} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3841};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3570, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3118} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4406} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3237} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3647};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4161, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3715} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3570} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4729} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5143};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4348 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3172 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4069 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4265, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3817} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4348} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4069};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4633 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3742 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3461 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3361, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4986} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3742} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4633} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3461};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3789 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4964 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4676 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3101, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4716} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4964} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3789} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4676};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4071, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3622} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3361} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4265} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3101};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4026 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4916 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3130 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4535, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4080} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4916} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4026} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3130};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 = !b_man[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4868 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934 = !a_man[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3201 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3695 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4792, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4342} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3201} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4868} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3695};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3410 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4587 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4302 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3631, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3177} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4587} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3410} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4302};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3167, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4784} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4535} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4792} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3631};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4139, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3688} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3167} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4071} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3309};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4474, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4020} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4139} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4551} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3379};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5068, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4615} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3980} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4474} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4878};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3855, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3406} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4161} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3673} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5068};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3855} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3628} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4532};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3786 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4514 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3623 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3334 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5075, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4621} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3623} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3334} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4514};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5079 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4793 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3900 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4168, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3719} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4793} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5079} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3900};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5123 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4231 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891 = !a_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3946 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3904, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3457} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4231} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5123} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3946};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4502, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4055} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4168} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5075} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3904};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 = !b_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5042 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 = !b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3865 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3494, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5106} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5042} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3865};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3874 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4766 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4344, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3896} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3874} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4766};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3582 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4757 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4479 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4394, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3937} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4757} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3582} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4479};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4462, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4011} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3896} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3494} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4394};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3629 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3911 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4803 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4129, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3679} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3911} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3629} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4803};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4190 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5087 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3294 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3224, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4842} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5087} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4190} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3294};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3333, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4953} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4842} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3679} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3937};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4833, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4383} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4011} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4502} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3333};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3287 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4468 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4181 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3265, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4885} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4468} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3287} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4181};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3374, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4999} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4621} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3719} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4885};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4748 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3857 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3573 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4435, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3987} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3857} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4748} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3573};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3600, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3144} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4435} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5106} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3265};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3977, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3527} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3374} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4055} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3144};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4165 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3269 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5061 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4894, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4447} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3269} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4165} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5061};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4451 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4727 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3554 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3995, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3540} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4727} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4451} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3554};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4774 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3882 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3604 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3731, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3272} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3882} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4774} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3604};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4585, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4136} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3995} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4894} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3731};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3235 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4130 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4481, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4028} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3235} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4130};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4405 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3227 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4251, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3807} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4405} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3227};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5016 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4122 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3838 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3089, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4704} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4122} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5016} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3838};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3686, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3232} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4251} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4028} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3089};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4281, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3831} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3457} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4585} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3686};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3957 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5131 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4847 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3860, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3413} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5131} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3957} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4847};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3343 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4522 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4241 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5034, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4575} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4522} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3343} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4241};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346 = !a_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4838 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4138 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5035 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3535, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3079} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5035} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4138};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4804, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4357} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4481} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4838} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3079};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4237, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3788} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4575} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3413} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4804};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4877, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4425} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4281} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4953} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3788};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3403, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5024} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3977} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4383} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4877};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3873 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5052 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4765 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4411, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3956} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5052} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3873} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4765};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3261 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4443 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4156 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3513, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5122} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3261} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4156};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4367, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3914} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3513} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4411} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4704};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3216 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4111 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5005 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3776, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3312} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4111} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5005};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4718 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3829 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3547 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4671, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4220} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3829} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4718} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3547};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3465, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5083} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3776} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3807} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4671};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3198, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4813} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3540} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4447} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3272};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3153, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4773} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3465} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4367} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3198};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3313 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4497 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3505 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4396 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4940, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4490} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3505} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4396};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4629, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4174} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4497} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4940};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3847 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5026 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4736 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3302, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4930} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5026} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3847} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4736};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4458 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3563 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3277 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4210, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3765} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3563} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4458} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3277};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3422, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5041} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4930} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4629} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3765};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4061, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3611} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4136} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3232} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5041};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4921, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4470} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3831} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3153} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4061};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4612, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4159} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3527} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4425} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4921};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3286, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4908} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4129} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3224} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5034};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4488 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3303 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3592 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3182, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4796} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3303} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4488} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3592};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4569 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3680 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4764, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4314} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3680} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4569} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3535};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4194, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3747} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4796} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3860} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4764};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3671, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3214} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4908} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4237} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3747};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5069 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4173 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3891 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5113, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4661} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4173} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5069} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3891};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3644, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3190} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3302} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5113} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4210};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3614 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4782 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4505 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3945, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3504} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4782} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3614} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4505};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4216 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3322 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5114 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4850, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4404} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3322} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5114};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4548, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4093} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4850} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3945} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3987};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5138, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4689} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4314} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4548};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4811 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3639 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4534 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4988, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4539} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4811} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4534};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5094 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4199 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3920 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4085, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3633} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4199} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5094} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3920};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4248 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5141 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3352 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3823, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3365} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5141} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4248} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3352};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5098, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4644} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3633} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4539} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3365};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3399 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4576 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4295 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3553, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3107} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4576} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3399} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4295};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4858 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3687 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3967 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4721, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4266} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3687} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4858} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3967};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3929, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3484} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4266} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3107} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3600};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4568, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4120} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5138} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3484};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3115, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4726} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4357} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3422} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3190};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4322, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3870} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3504} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4404};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4018, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3566} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4093} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4322} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4999};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3710, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3257} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3115} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4689} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4018};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4304, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3853} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4120} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3214} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3710};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4612} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5024} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3853};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3888, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3437} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3823} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4721} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3553};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5054, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4603} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3182} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4085} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4988};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3355, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4979} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4603} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3437} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4194};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4000, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3546} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3671} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4979} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4568};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3082 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3979 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4255 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3518, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5127} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3979} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3082} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4255};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3694 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4871 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4586 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4416, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3966} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3694} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4586} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4871};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4305 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3409 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3129 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3248, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4866} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3409} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4305} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3129};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3625, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3171} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3966} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5127} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4866};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4025 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3601 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4775 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4046, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3590} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3601} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4775};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4149, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3699} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4025} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4344} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3590};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4529, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4074} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4462} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3286} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3699};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3096, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4710} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3171} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4833} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4074};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3314 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4498 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4208 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4944, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4494} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4498} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3314} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4208};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3930 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5104 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4822 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3779, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3321} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5104} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3930} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4822};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4545 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3649 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3362 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4679, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4225} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3649} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4545} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3362};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4786, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4334} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3321} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4494} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4225};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4257, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3813} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5098} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3929} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4334};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4900, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4452} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3813} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4710} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3403};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4304} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3546} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4452};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4487, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4034} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3518} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4679} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4416};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3612 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4506 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4634, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4180} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3612} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4506};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3581, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3128} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4944} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4180} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3779};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4856, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4408} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3625} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4034} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3128};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4553 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3372 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4263 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3205, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4821} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3372} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4553} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4263};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3988 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3091 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4880 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4109, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3661} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3091} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3988} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4880};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4595 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3703 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3419 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5014, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4563} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3703} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4595} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3419};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4215, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3772} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4821} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4563};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4217 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3323 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5111 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3472, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5088} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3323} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5111};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3659 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3938 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4829 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4373, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3922} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4829} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3659} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3938};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3311, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4937} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5088} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3248} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3922};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3691, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3239} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4937} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3772} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4529};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3426, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5046} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4257} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3239};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3137 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4315 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4035 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3846, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3393} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4315} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3137} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4035};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5119, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4670} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3393} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4149} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5054};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4926 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3754 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4744, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4298} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3754} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4926} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4046};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3955, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3510} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4298} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3888} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4786};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4592, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4140} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4670} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3355} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3510};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4327, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3877} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3096} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4140} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4000};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5046} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4900} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3877};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3947 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4228 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5120 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4969, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4519} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4228} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3947} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5120};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4810, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4363} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5014} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3846} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4519};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4839 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3668 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4561 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3804, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3347} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3668} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4839} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4561};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4275 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3100 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3384 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4702, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4249} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3100} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4275} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3384};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3650, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3195} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4249} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4744};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3121, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4733} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4215} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3195};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3761, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3300} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3691} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4733} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4592};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4649 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3762 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3477 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4172, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3728} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3762} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4649} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3477};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3383, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5004} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3728} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3581} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4487};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3912, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3463} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3205} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4109} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4373};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4515 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3335 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4065, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3616} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3335};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5080, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4625} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4634} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3616} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3472};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4287, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3836} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4625} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3463} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3311};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4928, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4478} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5004} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4856} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3836};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3430 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4323 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4604 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4444, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3991} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4323} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3430} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4604};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4890 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3996 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3714 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3538, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3086} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3996} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4890} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3714};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4042 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4938 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3145 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3270, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4892} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4042} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4938} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3145};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4554, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4099} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3086} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3991} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4892};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4024, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3571} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5119} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4099} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3955};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4658, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4207} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3571} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4478} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3426};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3300} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4327} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4207};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3344 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5132 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3958 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3229, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4846} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5132} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3344} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3958};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4570 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3677 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4848 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4134, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3683} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3677} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4570} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4848};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3982, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4846} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3683};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4898 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4008 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3724 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3868, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3417} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4008} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4898} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3724};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3112 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3394 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4285 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5038, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4582} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3112} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3394} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4285};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3441 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4613 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4330 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4769, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4319} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4613} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3441} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4330};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4882, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4433} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4582} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3417} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4319};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4352, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3901} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4554} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3532} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4433};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4659 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3773 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3489 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4510, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4058} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3773} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4659} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3489};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4051 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3154 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4945 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3607, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3152} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3154} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4051} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4945};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3717, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3152} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4058} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3912};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3186, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4802} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3262} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3383} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4287};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4995, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4546} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4024} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3901} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4802};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4380 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3468 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4238 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4401, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3944} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3468} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4238};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3339, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4959} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4380} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4065} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3944};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4617, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4164} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4810} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5080} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4959};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4242, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3795} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4702} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3804} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4969};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5145, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4693} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3270} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4444} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3538};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3452, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5070} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3795} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3650} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4693};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4089, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3640} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4164} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3121} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5070};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3828, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3370} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4928} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3640} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3761};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4546} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4658} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3370};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22954 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4664 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3496 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4456, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4005} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4664} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3496};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3767 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4655 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4870, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4419} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3767} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4655};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4374 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3486 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3196 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3702, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3251} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3486} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4374} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3196};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4823, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4377} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4870} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4005} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3702};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3878, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3429} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5122} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3956} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4823};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3533 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4701 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4422 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3440, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5057} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4701} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3533} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4422};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4989 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4094 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3811 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4606, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4154} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4094} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4989} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3811};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3206 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4385 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4102 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3281, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4902} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4385} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4102};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3665, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3208} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4606} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3440} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4902};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3539 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3252 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4432 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5091, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4638} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3252} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3539} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4432};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4137 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3242 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3757 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4932 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4121, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3674} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3757} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4932};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4337, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3890} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3242} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4137} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4121};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3819 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11781 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4709 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4182, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3741} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11781} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3819} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4709};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4565, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4110} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4337} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3741};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4300, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3849} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3208} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4377} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4110};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3595 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3240, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4861} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3595} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4456} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4490};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4143, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3693} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4182} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5091} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3281};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4781, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4329} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3665} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4861} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3693};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4521, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4068} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4300} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4329};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4101, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3654} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3240} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4143};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3840, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3386} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4813} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3878} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3654};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5044 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4145 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3864 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3925, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3474} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4145} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5044} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3864};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5050, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4594} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3925} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3312} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4220};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5007, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4556} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5083} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5050} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3914};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4645 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3475 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4365 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5028, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4573} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3475} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4645} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4365};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4082 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3188 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4980 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3856, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3405} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3188} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4082} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4980};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3175, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4790} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4419} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5028} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3856};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4692 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3803 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3523 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4756, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4308} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3803} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4692} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3523};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4078, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3627} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3251} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4756} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4154};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3396, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5018} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3474} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3175} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4078};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3619, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3164} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4565} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4594} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3396};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4734, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4290} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4781} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4556} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3619};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3386} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4521} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4290};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4963, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4511} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3870} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4101} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5007};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3796, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3342} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4773} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3840};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4511} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4734} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3342};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3756, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3293} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4726} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4963};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3796} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4470} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3293};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3257} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3756} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4159};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22921 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3325, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4949} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3405} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4308} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4573};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3816, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3360} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3890} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3325} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4790};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4031 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4923 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4271, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3826} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4031} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4923};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4414 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3594, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3141} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4414} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4271} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3674};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3794 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4970 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4683 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4913, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4466} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4970} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3794} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4683};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3179 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4354 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4073 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4015, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3558} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4354} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3179} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4073};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4636 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3748 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3466 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3111, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4723} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3748} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4636} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3466};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4496, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4048} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4015} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4913} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3111};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4981, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4533} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5057} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3594} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4496};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3132, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4747} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4981} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3816} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5018};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3164} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3132} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4068};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3124 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4022 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3259, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4879} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3124} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4022};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4335 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4619 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3444 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4957, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4504} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3444} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4335} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4619};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4903 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4013 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3729 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4057, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3603} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4013} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4903} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3729};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4800, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4347} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4957} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4879} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4057};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3485, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5101} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3558} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4466} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4800};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4345 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3458 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3168 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5067, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4616} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3458} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4345} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3168};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4960 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4064 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4292 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3117 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3148, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4768} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4292} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3117};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3899, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3450} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4064} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4960} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3148};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4647, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4195} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3899} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5067} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4723};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5130, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4682} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4647} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3485} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4949};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3738 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4914 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4627 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4162, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3713} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4914} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3738} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4627};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3750, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3289} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3259} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3826} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4162};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4230, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3783} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3750} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3141} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4048};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4713, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4259} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3627} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4533} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4230};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3360} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5130} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4259};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3849} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4713} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4747};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22578 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3160 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3389 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4283 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3941, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3499} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3389} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4283};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3791, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3338} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3941} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3160} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4768};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3636, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3185} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3713} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4616} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3791};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4387, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3934} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3289} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3636} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4195};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4387} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3783} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4682};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4609 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3720 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3435 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3682, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3226} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3720} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4609} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3435};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4003 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3108 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4895 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4844, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4398} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3108} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4003} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4895};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4691, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4240} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4844} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3682} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3603};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4544, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4087} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3450} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4691} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4347};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5101} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4544} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3934};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4558 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3378 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3568, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3119} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4558} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3378};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3097 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4272 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3993 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4475, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4021} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4272} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3097} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3993};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4579, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4132} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3568} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4475};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3530, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5140} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4504} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3338};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3530} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3185} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4087};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4477 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4260 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3367 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3087 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5000, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4552} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3367} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4260} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3087};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3358 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4541 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4252 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11794 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4358, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3910} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4541} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3358} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4252};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3917 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4807 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3723, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3917} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4807};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4817 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3646 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3460, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5076} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4817} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3646};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3194, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5076} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3723} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3910};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4358} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4552} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3194};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3711 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4886 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3656 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4550 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4097, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3645} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3656} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4550};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3297, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4925} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4886} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3711} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4097};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3985 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3834, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3985} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3460} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3645};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4206, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3759} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3119} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5000} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4021};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3834} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4925} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3759};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3700 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4531 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3637 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5084 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3907 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4889, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5084} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3907};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3637} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4531} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4889};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4680 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4798 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4440);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3268 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4171);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4226 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4680)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4226);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4624 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4809);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3380 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4282);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3249 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3700)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3249);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4730 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4654);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3416, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5037} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4398} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3226} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3297};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4132} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5037};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4530 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5108 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3863);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4075 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4530) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4075);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3416} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4240} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5140};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3737 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4317 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3981);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4428 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4992);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3279 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3737 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3279);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3369 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4834);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3218 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3522);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4027 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4477)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4027);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3970 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3099);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3548 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3585);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4038 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4972);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22570 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22578)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22570);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3351 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5045 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5045;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3575 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4246);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4697 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4202);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4652 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5064);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3447 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4755);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4516 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22911 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4968)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4516);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22921) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22911);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3136 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3278);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3736 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22743);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22737 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22737;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22749 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22757);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22731 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22739);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22745 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22922 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22745;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22934 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22951 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22922);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22954)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4402 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11813 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3222 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4007, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3552} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11813} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4402} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3222};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4976, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4525} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4007} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4675};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3810, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3354} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3244} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4413} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4147};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5043, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4591} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4976} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4212} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3810};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4371 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4891;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3968 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3562, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3113} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4371} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3968};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4113 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5142 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3090;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3684 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4737 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3133);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4859 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3655 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4467, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4016} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3684} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5142} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4859};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4907, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4457} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4113} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3562} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4467};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4707, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4254} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5051} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3884} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4907};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3875, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3424} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5115} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4707} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3953};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3296, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4924} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3875} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5043} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4284};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4954 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3448 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3780 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4990 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4667 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4463 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4845);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4836, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4390} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3780} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4954} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4667};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4059 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3978 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3260);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3162 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4801 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4955);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4338 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3861 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4273);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3936, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3491} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3162} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4059} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4338};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4391 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3500 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3299 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3931);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3211 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3675, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3221} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3500} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4391} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3211};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4639, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4188} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3936} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4836} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3675};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4017 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3120 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3176 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4905 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3906 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4232);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4198, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3753} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3120} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4017} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4905};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4622 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4922 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3732 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4758 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3376);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3451 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4395 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3751);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5102, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4648} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3732} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4622} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3451};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4577 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3666 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3766);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3400 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4184 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4851);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4296 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4324 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4715);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3291, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4917} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3400} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4577} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4296};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3743, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3283} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5102} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4198} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3291};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3480, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5092} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4342} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4080} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3177};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3543, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3093} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3743} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3480};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4379, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3927} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4716} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3817} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4986};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4450, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3998} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3622} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4784} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4379};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4777, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4325} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3543} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4853} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4450};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4205, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3758} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3118} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4777} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4020};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3898, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3449} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3296} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3715} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4205};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4572} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3898} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3406};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4574, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4126} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4401} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3113} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3229};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3407, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5030} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5038} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4134} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3868};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3210, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4828} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3552} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4574} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3407};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3276, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4897} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4525} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3354};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3613, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3159} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3688} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4591} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3276};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4311, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3858} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4510} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3607} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4769};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3142, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4761} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4016} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3753} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4917};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4115, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3667} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4457} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4311} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3142};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4049, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3596} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4390} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4648} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3491};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5020, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4566} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3283} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4049} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4188};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4177, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3734} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4254} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4115} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5020};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4517, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4062} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4177} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3424} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4325};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5107, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4657} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3613} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4924} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4517};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4615} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5107} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3449};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4950, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4500} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3221} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3339} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4242};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3850, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3398} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5092} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4950} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3927};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5086, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4632} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3850} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3093} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3998};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3785, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3327} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4126} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5145} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5030};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4684, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4233} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3982} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3858} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4882};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4752, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4301} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3785} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4828} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4684};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3918, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3471} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4752} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4897} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3734};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3345, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4966} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5086} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3159} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3918};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3758} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3345} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4657};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3524, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5134} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3717} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4761} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3596};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3586, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3134} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3667} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3524};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4421, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3972} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4500} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4617} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3452};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4492, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4041} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4421} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3398} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4301};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4819, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4370} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3586} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4632} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4492};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4062} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4819} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4966};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4155, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3706} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3186} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5134} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3972};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3253, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4872} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3327} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4233} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4352};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5060, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4608} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4089} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4872} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4995};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3706} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3828} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4608};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3318, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4941} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3253} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3134} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4155};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4041} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5060} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4941};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3471} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3318} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4370};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22928 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4725 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3442);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3892 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3777);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3192 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3192;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4221 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3200);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3658 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3802);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5002 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22938 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5002;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22933) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22938);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4247 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3498);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3943 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4350);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4732 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4732;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4799 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4307);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4759 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3359);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4473 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22919 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4473;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22947 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22931) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22919);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22917 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22958)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22947);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22928 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22917);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3815 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3584);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4039 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4974);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3350 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3388);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3839 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5040);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3942 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4399)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3942);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3421 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3722);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4167 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3565);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4019 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4578);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5033 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4688);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4958 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4430 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3336)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4958);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4881) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4430);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5139 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3895);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4346 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4270);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4720 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3746);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4382 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4193);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3897 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5032 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4349)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3897));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3427 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3408)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5032);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3328 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3427;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3786)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3328);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3818 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3404;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3801 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4672;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4708 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3670, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3215} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3801} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3818} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4708};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5097} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3215} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3932};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4119 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4832);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3544 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4946;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4700 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4144;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4700} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3544} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3670};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5023 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4571);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3975) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[45] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4407);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3487 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3952 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3236) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4852);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4002 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3652 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3487) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4002);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[45] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[45]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4032 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3577));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3837 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3837);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4151 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3135 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4288 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3516 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3135 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3531);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4601 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4127 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3516;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4050 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3866;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3598 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3414;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4050)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3598);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[39] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4601) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4151);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4412)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3959);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3411 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[40] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3411;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[40]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[39]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3126 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4742));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3149;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4867 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3588 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3572 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3605));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3246 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4840 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3588;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[38] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3246) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4867);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[39]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[38]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4293 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3844));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3964 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3520 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3492) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[37] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3520) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3964);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[38]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[37]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4200 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3391 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5010));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[36] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4200) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3916;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[37]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[36]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7499 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4788 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4523 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5110 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3169 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4053 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4523;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[42] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3169) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4788);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3506 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5117));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4665;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4223 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4614);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3301 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4211;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4163) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3763)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3301);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4448 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4223 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4448;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3331) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4542;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[43] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[43]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[42]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[44] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22802) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[43]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7493 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[44];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4560 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4106));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4116 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4364 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4812)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4364);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4641 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4116 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4677 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4641;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4227 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4919) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4580;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[35] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4227) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4677);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[36]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[35]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3657 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3203));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4204;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4717 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4656));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3319 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4717;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4947 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3564) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4100;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[34] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4947) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3319);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[35]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11804) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[34]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4818 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4369));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3591 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4044 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4279) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[33] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4044) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3591);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[34]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[33]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4997 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3919 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3470));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[32] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4218 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4997;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[33]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[32]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7532 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4166;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4825 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454);
assign N11217 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22915;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006 = !N11217;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4918 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3718;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4375 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3292)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4918);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4825) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4375);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4355 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[30] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4355;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5085 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4631));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4306 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4179) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4753 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3733) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3642;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4753) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3315) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4306);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[31]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[30]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[32]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[31]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3275 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4899));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5025 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3402 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5073;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5103 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4454;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4651 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4006;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5103) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4651);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[29] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3402) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5025);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[30]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[29]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3721 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4449 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3997));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[28] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4491 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3721;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[29]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11803) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[28]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7433 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7532 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7433);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3770 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3308));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3886 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4485;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3438 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4762) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4933;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[41] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3438) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4815) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3886);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[42]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[41]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[41]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[40]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7505 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7499) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7493) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3545 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3092));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3672 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4118 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4438;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4694) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4244);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[27] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4118) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3672);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[28]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[27]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3080 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4706 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4256));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[26] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3583 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3080;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[27]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[26]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3809 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3353));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4831 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4384 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11836 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4261;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11836;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4384) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4831);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[26]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[25]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4512 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4978 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4524));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[24] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4837) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4512;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[25]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[24]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7467 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22759 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3624));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5096 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3482 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3155;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4091 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3151;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3434 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4091 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3434 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4771);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[23] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3482) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5096);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[24]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[23]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7467 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7429 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7505 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3871 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3166 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4783));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[22] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3871 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4392;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22612 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[23]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11805) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663 = !rm[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679 = !rm[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22613 = !((rm[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788 = (!a_sign) ^ b_sign;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666 = !rm[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684 = !((rm[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5 = (rm[0] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22637 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22613 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22622 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7679 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7663) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4862 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4415));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3821 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4269 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3305;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3418;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[17] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4269) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3821);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3455 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3556 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3455;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3105 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4662) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3349;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[18] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3105) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3556);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[18] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[18]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[17]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4029 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3962 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3514));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[16] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4029;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[17] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[17]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[16]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7731 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[18] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[17]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22569 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22566 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22575));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22579 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22563 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22579);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22569) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22563;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22560 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5126 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4674));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[15] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3778) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22560;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[15] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[15]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47]) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[14]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[16] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[16]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[15]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7742 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[15] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[16]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7751 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7731 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7742);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3479 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4336 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3887));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[13] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4092 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3479;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[14] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[14]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[13]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4187 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3436 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5056));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3606) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4187;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[13] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[13]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[12]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7753 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[14] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[13]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4874 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4857 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4874 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4906 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4602 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4148));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[11] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4857 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4906;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[12] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[12]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[11]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3551 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3701 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3247));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[10] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4286 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3551;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[11] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[11]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11801) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[10]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7763 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[12] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[11]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7761 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7753 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7763);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22628 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7761 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5077) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4178;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5136 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4754 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4303));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3854) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5136;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[2]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47]) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[0] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3346 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3620;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[0] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[0] | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[1] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[1]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[0]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7749 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7729 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7749);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4333 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3883));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3745 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4192 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4588;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[21] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4192) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3745);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[22] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[22]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[21]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3233 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3431 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5053));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[20] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5058 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3233;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[21] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[21]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[20]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7759 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[22] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[21]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4599 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4146));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3698;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5093 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3158);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3618 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3243;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4776) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4066)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3618);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3373 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5093 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4911 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3373;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4460 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3949) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3083;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[19] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4460) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4353) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4911);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[20] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[20]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[19]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[19] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[19]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11802) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[18]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7721 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[20] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[19]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7740 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7759 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7721);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7744 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7729 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7740);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3385 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4264 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4865 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4418));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[9] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3385 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4264;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[10] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[10]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[9]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4985 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3965 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3517));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4971) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4985;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[9] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[9]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[8]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7725 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[10] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3630 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5129 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4678));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[7] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3954 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3630;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[8] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[8]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[7]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4341 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4224 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3782));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4746) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4341;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[7] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[7]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[6]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7735 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7723 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7725 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7735);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4423 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3589 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3139));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4528 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4423;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[3] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[3]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[2]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3708 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4495 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4045));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3999) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3708;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[4] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[4]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[3]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7757 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[3] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5062 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3320 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4943));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[5] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3473 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N5062;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[6] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[6]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[5]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[5] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[5]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11800) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[4]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7746 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[6] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7733 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7757 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7746);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7738 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7723 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7733);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22638 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7744 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7738;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22628 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22638);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22619 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22615 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22622 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22619);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22614 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22637 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22615);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22617 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22646;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22631 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22643 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22634);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22641 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22617 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22631);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22614) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22612)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22641);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8524 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8524;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11903 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7429 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8421 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[45] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11903;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3008 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3012 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3008 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3012);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2885 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2889 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2885 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2889);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__7 = (rm[0] & rm[1]) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7666;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8254 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__7) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7684) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__5) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8254);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2919 = !(a_exp[7] & a_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2917 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11829 = !((a_exp[0] & a_exp[1]) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2917);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2919 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11829);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2955 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2959 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2934) | a_man[0]) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2955) | a_man[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2940 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2961 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2950 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2971 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2953 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2940 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2961) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2950) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2971);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2965 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2975 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2959) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2953) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2965) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2975);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2796 = !(b_exp[7] & b_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2794 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11821 = !((b_exp[0] & b_exp[1]) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2794);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2796 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11821);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2832 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2836 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2811) | b_man[0]) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2832) | b_man[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2817 = !(b_man[10] | b_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2838 = !(b_man[6] | b_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2827 = !(b_man[8] | b_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2848 = !(b_man[4] | b_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2830 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2817 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2838) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2827) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2848);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2842 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2852 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2836) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2830) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2842) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N2852);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__19 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__17));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__12 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__10));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3051 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__13) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3051) | (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__20 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__14 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__21;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8319 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857 = !a_exp[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888 = !(b_exp[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7890 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852 = !(a_exp[6] & b_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897 = !(a_exp[5] & b_exp[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861 = !(a_exp[4] & b_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908 = !(a_exp[3] & b_exp[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7865 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870 = !(a_exp[2] & b_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916 = !(a_exp[1] & b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7903 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879 = b_exp[0] | a_exp[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900 = !(a_exp[1] | b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854 = !(a_exp[2] | b_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7885 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7903)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7885);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892 = !(a_exp[3] | b_exp[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920 = !(a_exp[4] | b_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881 = !(a_exp[5] | b_exp[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913 = !(a_exp[6] | b_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7863 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7849 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7882)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7863);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7865) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7849);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867 = !(b_exp[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7869 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9] = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7890)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7869);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7915 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7899 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7857) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7899) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7915);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7868 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7888 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7867));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7868;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8228 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8228;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8319 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8507 = b_man[21] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8511 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[21]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8507);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8545 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8545;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8467 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8511) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7852 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7913));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7864 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7923 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7898) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7907 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7894;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7891 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7873;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7907) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7891);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[6] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7923) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7864));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8015 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7870 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7854));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7918 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7904 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7848) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7904) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7918));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7878 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7916 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7900));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7879) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7878;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684 = !b_exp[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696 = !a_exp[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0] | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7902 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7902;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7881 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7897));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7861 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7920));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7874 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7892;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7895 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7871) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7908;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[4] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7895) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7859) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7874));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11840 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11840);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8015) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3109;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3390 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3560));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3095 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3390;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4711 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3690) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4584;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[46] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N4711) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3095);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[47] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[46] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11807));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[46] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[46]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[45]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22795) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22815 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22806) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3973) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22798));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22788 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22815) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22804 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22810) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22819) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22816));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22792 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22818) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11806) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22804));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22788 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22792);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7506 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[47] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[46]) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7540 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7534 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7506 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7540);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7473 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7469 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7486 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7469 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7486;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7473 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7511 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7511 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[24] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7534 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[24]) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[47]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[8]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8018 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8018) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[7] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[7]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7991));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[6] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[6]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8004));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8136 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22677 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684 & a_exp[0]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22684) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22696));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[0] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22677;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[1]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8132 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[0] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8130 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8136 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8132);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22861 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22856 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22861) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22871 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22852) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22869 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22848) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7875) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22875));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7998);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22865 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22869) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22872 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22865) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22871));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8140 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22856 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22872);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[2] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8014 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[2]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8047 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7994 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[3]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8047);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8127 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8134 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8140 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8127);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8138 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8130 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8134);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7990 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7993 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8011);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8016 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7990 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8001);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8016;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[9]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[9]);
assign N11222 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8157 = !N11222;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22706 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8138 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[8]) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8157);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22861) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22846);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8176 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[8]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22987 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22854 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[5] = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[5] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22987;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8181 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[5] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1861);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8187 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8176 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8181);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8178 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8188 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8173 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6] | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8190 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8188 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8173);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8183 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8178 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8190);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8206 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8212 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8206 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22693 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8212) | (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8187 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8183);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22685 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22706 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22693);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__49 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22685;
assign x[21] = !((N11181 & N10691) | ((!N11181) & N10693));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7473 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7511;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7484 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7540 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7441) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7551 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7484);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11896 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7551 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8374 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[44] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11896;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8411 = b_man[20] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8463 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[20]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8411);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8420 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8463) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[20] = !((N11175 & N10698) | ((!N11175) & N10700));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7479 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7513 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7527);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7517 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7545 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7430);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7530 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7516 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7530;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7447 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7463);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7478 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7497);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7446 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7462 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7517) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7479)) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7446);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7462;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8547 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[19]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[43]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8536 = b_man[19] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8415 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[19]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8536);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8371 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8415) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[19] = !((N11178 & N10705) | ((!N11178) & N10707));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7521 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7538;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7424 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7440;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7520 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7452 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7469;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7481 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7486 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7504;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7512 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7520) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7481) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[18] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7512) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8497 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[18]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[42]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8442 = b_man[18] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8368 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[18]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8442);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8543 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8368) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[18] = !((N11176 & N10712) | ((!N11176) & N10714));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7433 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7467);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7422 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7532) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7499)) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[17] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7422;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8452 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[17]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[41]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8342 = b_man[17] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8539 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[17]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8342);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8494 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8539) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[17] = !((N11177 & N10719) | ((!N11177) & N10721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7439 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7468 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11889 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7439 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8403 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[40] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11889;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8468 = b_man[16] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8489 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[16]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8468);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8450 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8489) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[16] = !((N11176 & N10726) | ((!N11176) & N10728));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7543 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7517 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7550);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7450 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7530);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7459 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7543 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[15] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7459) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8352 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[15]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[39]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8373 = b_man[15] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8446 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[15]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8373);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8400 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8446) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[15] = !((N11180 & N10733) | ((!N11180) & N10735));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7455 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7490);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7437 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7526 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7548);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7432 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7437;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7432) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8526 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[14]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[38]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8495 = b_man[14] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8396 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[14]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8495);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8351 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8396) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[14] = !((N11179 & N10740) | ((!N11179) & N10742));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7537 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7428 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7482);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[13] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7537) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8477 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[13]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[37]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8401 = b_man[13] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8346 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[13]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8401);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8522 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8346) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[13] = !((N11179 & N10747) | ((!N11179) & N10749));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7508 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7503 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7500);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7508) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8432 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[12]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[36]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8525 = b_man[12] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8519 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[12]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8525);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8474 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8519) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[12] = !((N11175 & N10754) | ((!N11175) & N10756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7476 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7446 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7476) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8383 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[11]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[35]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8430 = b_man[11] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8470 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[11]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8430);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8429 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8470) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[11] = !((N11178 & N10761) | ((!N11178) & N10763));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7491 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7520 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7443);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11882 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7491 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8556 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[34] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11882;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8554 = b_man[10] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8423 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[10]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8554);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8381 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8423) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[10] = !((N11177 & N10768) | ((!N11177) & N10770));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7475 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7461 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7475) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8506 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[9]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[33]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8458 = b_man[9] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8377 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[9]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8458);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8553 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8377) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[9] = !((N11178 & N10775) | ((!N11178) & N10777));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7495) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8459 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[8]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[32]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8361 = b_man[8] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8549 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[8]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8361);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8504 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8549) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[8] = !((N11175 & N10782) | ((!N11175) & N10784));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11875 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7524 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8410 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[31] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11875;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8484 = b_man[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8499 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[7]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8484);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8457 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8499) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[7] = !((N11180 & N10789) | ((!N11180) & N10791));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7437;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11868 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8363 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[30] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11868;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8390 = b_man[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8454 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[6]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8390);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8408 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8454) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[6] = !((N11180 & N10796) | ((!N11180) & N10798));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7464) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8535 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[5]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[29]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8512 = b_man[5] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8404 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[5]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8512);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8360 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8404) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[5] = !((N11180 & N10803) | ((!N11180) & N10805));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7436) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8486 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[4]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[28]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8417 = b_man[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8354 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[4]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8417);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8533 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8354) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[4] = !((N11175 & N10810) | ((!N11175) & N10812));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11861 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7470 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8440 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[27] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11861;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8541 = b_man[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8529 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[3]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8541);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8483 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8529) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[3] = !((N11178 & N10817) | ((!N11178) & N10819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11854 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7481 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8391 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[26] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11854;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8447 = b_man[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8479 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[2]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8447);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8439 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8479) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[2] = !((N11177 & N10824) | ((!N11177) & N10826));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11847 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7546 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8341 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[25] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11847;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8348 = b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8434 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[1]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8348);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8388 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8434) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[1] = !((N11177 & N10831) | ((!N11177) & N10833));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8515 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[0]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8347) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[24]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8472 = b_man[0] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8384 = (float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_man[0]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8472);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8337 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8384) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8416) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47));
assign x[0] = !((N11176 & N10838) | ((!N11176) & N10840));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7522 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7419 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7435;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7456 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7485) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7522) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7494) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7425);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N7456) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[46];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8324 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[22]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__44) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[46]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8329 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__47 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26);
assign x[22] = !((N11175 & N10894) | ((!N11175) & N10896));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469 = float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__32;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8288 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26);
assign x[30] = !((N11179 & N10852) | ((!N11179) & N10847));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8282 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[6];
assign x[29] = !((N11179 & N10852) | ((!N11179) & N10854));
assign x[28] = !((N11179 & N10852) | ((!N11179) & N10861));
assign x[27] = !((N11176 & N10852) | ((!N11176) & N10868));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8263 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[3];
assign x[26] = !((N11177 & N10852) | ((!N11177) & N10875));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8285 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N1054;
assign x[25] = !((N11176 & N10852) | ((!N11176) & N10882));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N8279 = !float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[1];
assign x[24] = !((N11178 & N10852) | ((!N11178) & N10889));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22682 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0] & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__38) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[0]) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22681));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22689 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N469 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__42));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22678 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N22689 | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__27) | float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26);
assign x[23] = !((N11180 & N10901) | ((!N11180) & N10903));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3068 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__22 & (!b_sign));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3074 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15 & a_sign) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3068));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[31] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N3074) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__26) & float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_N11788));
reg x_reg_31__I2040_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I2040_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[31];
	end
assign x[31] = x_reg_31__I2040_QOUT;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__24[44] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__25[23] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__30[0] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[4] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__31[5] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[1] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[2] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[3] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[6] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[7] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[10] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[16] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[20] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[21] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__45[23] = 1'B0;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_0_inst_inst_cellmath__48[2] = 1'B0;
endmodule

/* CADENCE  vLDwSgDWqxw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



