/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:20 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2876250654_bdw (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__10,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23;
wire [47:0] inst_cellmath__24,
	inst_cellmath__25;
wire  inst_cellmath__26,
	inst_cellmath__27,
	inst_cellmath__28;
wire [9:0] inst_cellmath__30,
	inst_cellmath__31;
wire  inst_cellmath__32,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42,
	inst_cellmath__44;
wire [24:0] inst_cellmath__45;
wire  inst_cellmath__46,
	inst_cellmath__47;
wire [9:0] inst_cellmath__48;
wire  inst_cellmath__49,
	inst_cellmath__51;
wire N440,N441,N442,N443,N444,N445,N446 
	,N447,N448,N449,N450,N461,N462,N463,N469 
	,N470;
cynw_cm_float_mul_ieee_inst_cellmath__17_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I0 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__19__2__bdw2876250654_bdw cynw_cm_float_mul_ieee_I1 (.inst_cellmath__19__2__out0(inst_cellmath__19), .inst_cellmath__19__2__in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__21_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I2 (.inst_cellmath__21_0_out0(inst_cellmath__21), .inst_cellmath__21_0_in0(inst_cellmath__19), .inst_cellmath__21_0_in1(inst_cellmath__17));
cynw_cm_float_mul_ieee_inst_cellmath__13__1__bdw2876250654_bdw cynw_cm_float_mul_ieee_I3 (.inst_cellmath__13__1__out0(inst_cellmath__13), .inst_cellmath__13__1__in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__26__9__bdw2876250654_bdw cynw_cm_float_mul_ieee_I4 (.inst_cellmath__26__9__out0({N441}), .inst_cellmath__26__9__in0(inst_cellmath__21), .inst_cellmath__26__9__in1(inst_cellmath__13));
cynw_cm_float_mul_ieee_inst_cellmath__10_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I5 (.inst_cellmath__10_0_out0(inst_cellmath__10), .inst_cellmath__10_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__12__0__bdw2876250654_bdw cynw_cm_float_mul_ieee_I6 (.inst_cellmath__12__0__out0(inst_cellmath__12), .inst_cellmath__12__0__in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__14_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I7 (.inst_cellmath__14_0_out0(inst_cellmath__14), .inst_cellmath__14_0_in0(inst_cellmath__12), .inst_cellmath__14_0_in1(inst_cellmath__10));
cynw_cm_float_mul_ieee_inst_cellmath__20__3__bdw2876250654_bdw cynw_cm_float_mul_ieee_I8 (.inst_cellmath__20__3__out0(inst_cellmath__20), .inst_cellmath__20__3__in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__26__8__bdw2876250654_bdw cynw_cm_float_mul_ieee_I9 (.inst_cellmath__26__8__out0({N440}), .inst_cellmath__26__8__in0(inst_cellmath__20), .inst_cellmath__26__8__in1(inst_cellmath__14));
cynw_cm_float_mul_ieee_inst_cellmath__15_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I10 (.inst_cellmath__15_0_out0(inst_cellmath__15), .inst_cellmath__15_0_in0(inst_cellmath__12), .inst_cellmath__15_0_in1(inst_cellmath__10));
cynw_cm_float_mul_ieee_inst_cellmath__22_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I11 (.inst_cellmath__22_0_out0(inst_cellmath__22), .inst_cellmath__22_0_in0(inst_cellmath__19), .inst_cellmath__22_0_in1(inst_cellmath__17));
cynw_cm_float_mul_ieee_inst_cellmath__26_1_bdw2876250654_bdw cynw_cm_float_mul_ieee_I12 (.inst_cellmath__26_1_out0(inst_cellmath__26), .inst_cellmath__26_1_in0({N441}), .inst_cellmath__26_1_in1({N440}), .inst_cellmath__26_1_in2(inst_cellmath__22), .inst_cellmath__26_1_in3(inst_cellmath__15));
cynw_cm_float_mul_ieee_inst_cellmath__23_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I13 (.inst_cellmath__23_0_out0(inst_cellmath__23), .inst_cellmath__23_0_in0(b_sign), .inst_cellmath__23_0_in1(a_sign));
cynw_cm_float_mul_ieee_inst_cellmath__41_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I14 (.inst_cellmath__41_0_out0(x[31]), .inst_cellmath__41_0_in0(inst_cellmath__26), .inst_cellmath__41_0_in1(inst_cellmath__23), .inst_cellmath__41_0_in2(inst_cellmath__22), .inst_cellmath__41_0_in3(inst_cellmath__15), .inst_cellmath__41_0_in4(b_sign), .inst_cellmath__41_0_in5(a_sign));
cynw_cm_float_mul_ieee_inst_cellmath__24_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I15 (.inst_cellmath__24_0_out0({inst_cellmath__24[47], inst_cellmath__24[46], inst_cellmath__24[45], inst_cellmath__24[44], inst_cellmath__24[43], inst_cellmath__24[42], inst_cellmath__24[41], inst_cellmath__24[40], inst_cellmath__24[39], inst_cellmath__24[38], inst_cellmath__24[37], inst_cellmath__24[36], inst_cellmath__24[35], inst_cellmath__24[34], inst_cellmath__24[33], inst_cellmath__24[32], inst_cellmath__24[31], inst_cellmath__24[30], inst_cellmath__24[29], inst_cellmath__24[28], inst_cellmath__24[27], inst_cellmath__24[26], inst_cellmath__24[25], inst_cellmath__24[24], inst_cellmath__24[23], inst_cellmath__24[22], inst_cellmath__24[21], inst_cellmath__24[20], inst_cellmath__24[19], inst_cellmath__24[18], inst_cellmath__24[17], inst_cellmath__24[16], inst_cellmath__24[15], inst_cellmath__24[14], inst_cellmath__24[13], inst_cellmath__24[12], inst_cellmath__24[11], inst_cellmath__24[10], inst_cellmath__24[9], inst_cellmath__24[8], inst_cellmath__24[7], inst_cellmath__24[6], inst_cellmath__24[5], inst_cellmath__24[4], inst_cellmath__24[3], inst_cellmath__24[2], inst_cellmath__24[1], inst_cellmath__24[0]}), .inst_cellmath__24_0_in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}), .inst_cellmath__24_0_in1({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__25_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I16 (.inst_cellmath__25_0_out0({inst_cellmath__25[47], inst_cellmath__25[46], inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24], inst_cellmath__25[23], inst_cellmath__25[22], inst_cellmath__25[21], inst_cellmath__25[20], inst_cellmath__25[19], inst_cellmath__25[18], inst_cellmath__25[17], inst_cellmath__25[16], inst_cellmath__25[15], inst_cellmath__25[14], inst_cellmath__25[13], inst_cellmath__25[12], inst_cellmath__25[11], inst_cellmath__25[10], inst_cellmath__25[9], inst_cellmath__25[8], inst_cellmath__25[7], inst_cellmath__25[6], inst_cellmath__25[5], inst_cellmath__25[4], inst_cellmath__25[3], inst_cellmath__25[2], inst_cellmath__25[1], inst_cellmath__25[0]}), .inst_cellmath__25_0_in0({inst_cellmath__24[47], inst_cellmath__24[46], inst_cellmath__24[45], inst_cellmath__24[44], inst_cellmath__24[43], inst_cellmath__24[42], inst_cellmath__24[41], inst_cellmath__24[40], inst_cellmath__24[39], inst_cellmath__24[38], inst_cellmath__24[37], inst_cellmath__24[36], inst_cellmath__24[35], inst_cellmath__24[34], inst_cellmath__24[33], inst_cellmath__24[32], inst_cellmath__24[31], inst_cellmath__24[30], inst_cellmath__24[29], inst_cellmath__24[28], inst_cellmath__24[27], inst_cellmath__24[26], inst_cellmath__24[25], inst_cellmath__24[24], inst_cellmath__24[23], inst_cellmath__24[22], inst_cellmath__24[21], inst_cellmath__24[20], inst_cellmath__24[19], inst_cellmath__24[18], inst_cellmath__24[17], inst_cellmath__24[16], inst_cellmath__24[15], inst_cellmath__24[14], inst_cellmath__24[13], inst_cellmath__24[12], inst_cellmath__24[11], inst_cellmath__24[10], inst_cellmath__24[9], inst_cellmath__24[8], inst_cellmath__24[7], inst_cellmath__24[6], inst_cellmath__24[5], inst_cellmath__24[4], inst_cellmath__24[3], inst_cellmath__24[2], inst_cellmath__24[1], inst_cellmath__24[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__45_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I17 (.inst_cellmath__45_0_out0({inst_cellmath__45[24], inst_cellmath__45[23], inst_cellmath__45[22], inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__45_0_in0({inst_cellmath__25[47], inst_cellmath__25[46], inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24]}));
cynw_cm_float_mul_ieee_inst_cellmath__5_1_bdw2876250654_bdw cynw_cm_float_mul_ieee_I18 (.inst_cellmath__5_1_out0(inst_cellmath__5), .inst_cellmath__5_1_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__31__bdw2876250654_bdw cynw_cm_float_mul_ieee_I19 (.inst_cellmath__44__31__out0({N446}), .inst_cellmath__44__31__in0(inst_cellmath__5), .inst_cellmath__44__31__in1(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__6_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I20 (.inst_cellmath__6_0_out0(inst_cellmath__6), .inst_cellmath__6_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__30__bdw2876250654_bdw cynw_cm_float_mul_ieee_I21 (.inst_cellmath__44__30__out0({N445}), .inst_cellmath__44__30__in0(inst_cellmath__6), .inst_cellmath__44__30__in1(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__8_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I22 (.inst_cellmath__8_0_out0(inst_cellmath__8), .inst_cellmath__8_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__4_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I23 (.inst_cellmath__4_0_out0(inst_cellmath__4), .inst_cellmath__4_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__34_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I24 (.inst_cellmath__34_0_out0(inst_cellmath__34), .inst_cellmath__34_0_in0({inst_cellmath__25[22], inst_cellmath__25[21], inst_cellmath__25[20], inst_cellmath__25[19], inst_cellmath__25[18], inst_cellmath__25[17], inst_cellmath__25[16], inst_cellmath__25[15], inst_cellmath__25[14], inst_cellmath__25[13], inst_cellmath__25[12], inst_cellmath__25[11], inst_cellmath__25[10], inst_cellmath__25[9], inst_cellmath__25[8], inst_cellmath__25[7], inst_cellmath__25[6], inst_cellmath__25[5], inst_cellmath__25[4], inst_cellmath__25[3], inst_cellmath__25[2], inst_cellmath__25[1], inst_cellmath__25[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__29__bdw2876250654_bdw cynw_cm_float_mul_ieee_I25 (.inst_cellmath__44__29__out0({N443}), .inst_cellmath__44__29__in0(inst_cellmath__34), .inst_cellmath__44__29__in1({inst_cellmath__25[24]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__28__bdw2876250654_bdw cynw_cm_float_mul_ieee_I26 (.inst_cellmath__44__28__out0({N444}), .inst_cellmath__44__28__in0({N443}), .inst_cellmath__44__28__in1(inst_cellmath__4));
cynw_cm_float_mul_ieee_inst_cellmath__44__27__bdw2876250654_bdw cynw_cm_float_mul_ieee_I27 (.inst_cellmath__44__27__out0({N447}), .inst_cellmath__44__27__in0(inst_cellmath__8), .inst_cellmath__44__27__in1({N446}), .inst_cellmath__44__27__in2({N445}), .inst_cellmath__44__27__in3({N444}));
cynw_cm_float_mul_ieee_inst_cellmath__44__26__bdw2876250654_bdw cynw_cm_float_mul_ieee_I28 (.inst_cellmath__44__26__out0({N448}), .inst_cellmath__44__26__in0({N447}), .inst_cellmath__44__26__in1({inst_cellmath__25[23]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__33__bdw2876250654_bdw cynw_cm_float_mul_ieee_I29 (.inst_cellmath__44__33__out0({N449}), .inst_cellmath__44__33__in0({N446}), .inst_cellmath__44__33__in1({N445}));
cynw_cm_float_mul_ieee_inst_cellmath__44__32__bdw2876250654_bdw cynw_cm_float_mul_ieee_I30 (.inst_cellmath__44__32__out0({N450}), .inst_cellmath__44__32__in0({N449}), .inst_cellmath__44__32__in1(inst_cellmath__34));
cynw_cm_float_mul_ieee_inst_cellmath__44_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I31 (.inst_cellmath__44_0_out0(inst_cellmath__44), .inst_cellmath__44_0_in0({N450}), .inst_cellmath__44_0_in1({N448}));
cynw_cm_float_mul_ieee_inst_cellmath__46_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I32 (.inst_cellmath__46_0_out0(inst_cellmath__46), .inst_cellmath__46_0_in0({inst_cellmath__45[24]}), .inst_cellmath__46_0_in1(inst_cellmath__44));
cynw_cm_float_mul_ieee_inst_cellmath__38_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I33 (.inst_cellmath__38_0_out0(inst_cellmath__38), .inst_cellmath__38_0_in0(inst_cellmath__46), .inst_cellmath__38_0_in1({inst_cellmath__24[47]}));
cynw_cm_float_mul_ieee_inst_cellmath__30_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I34 (.inst_cellmath__30_0_out0({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}), .inst_cellmath__30_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}), .inst_cellmath__30_0_in1({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__31_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I35 (.inst_cellmath__31_0_out0({inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}), .inst_cellmath__31_0_in0({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__48_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I36 (.inst_cellmath__48_0_out0({inst_cellmath__48[9], inst_cellmath__48[8], inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}), .inst_cellmath__48_0_in0(inst_cellmath__38), .inst_cellmath__48_0_in1({inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}), .inst_cellmath__48_0_in2({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__51__49__bdw2876250654_bdw cynw_cm_float_mul_ieee_I37 (.inst_cellmath__51__49__out0({N461}), .inst_cellmath__51__49__in0({inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__51__48__bdw2876250654_bdw cynw_cm_float_mul_ieee_I38 (.inst_cellmath__51__48__out0({N462}), .inst_cellmath__51__48__in0({N461}), .inst_cellmath__51__48__in1({inst_cellmath__48[8]}));
cynw_cm_float_mul_ieee_inst_cellmath__51_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I39 (.inst_cellmath__51_0_out0(inst_cellmath__51), .inst_cellmath__51_0_in0({N462}), .inst_cellmath__51_0_in1({inst_cellmath__48[9]}));
cynw_cm_float_mul_ieee_inst_cellmath__28_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I40 (.inst_cellmath__28_0_out0(inst_cellmath__28), .inst_cellmath__28_0_in0(inst_cellmath__20), .inst_cellmath__28_0_in1(inst_cellmath__13));
cynw_cm_float_mul_ieee_inst_cellmath__27_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I41 (.inst_cellmath__27_0_out0(inst_cellmath__27), .inst_cellmath__27_0_in0(inst_cellmath__21), .inst_cellmath__27_0_in1(inst_cellmath__14));
cynw_cm_float_mul_ieee_inst_cellmath__50__50__bdw2876250654_bdw cynw_cm_float_mul_ieee_I42 (.inst_cellmath__50__50__out0({N463}), .inst_cellmath__50__50__in0({inst_cellmath__48[9], inst_cellmath__48[8], inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__49_1_bdw2876250654_bdw cynw_cm_float_mul_ieee_I43 (.inst_cellmath__49_1_out0(inst_cellmath__49), .inst_cellmath__49_1_in0(inst_cellmath__51), .inst_cellmath__49_1_in1({N463}), .inst_cellmath__49_1_in2({inst_cellmath__48[9]}), .inst_cellmath__49_1_in3(inst_cellmath__28), .inst_cellmath__49_1_in4(inst_cellmath__27), .inst_cellmath__49_1_in5(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__37__43__bdw2876250654_bdw cynw_cm_float_mul_ieee_I44 (.inst_cellmath__37__43__out0({N470}), .inst_cellmath__37__43__in0(inst_cellmath__27), .inst_cellmath__37__43__in1(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__32__11__bdw2876250654_bdw cynw_cm_float_mul_ieee_I45 (.inst_cellmath__32__11__out0({N442}), .inst_cellmath__32__11__in0({inst_cellmath__30[8], inst_cellmath__30[7]}));
cynw_cm_float_mul_ieee_inst_cellmath__32__10__bdw2876250654_bdw cynw_cm_float_mul_ieee_I46 (.inst_cellmath__32__10__out0(inst_cellmath__32), .inst_cellmath__32__10__in0({N442}), .inst_cellmath__32__10__in1({inst_cellmath__30[9]}));
cynw_cm_float_mul_ieee_inst_cellmath__37__42__bdw2876250654_bdw cynw_cm_float_mul_ieee_I47 (.inst_cellmath__37__42__out0({N469}), .inst_cellmath__37__42__in0(inst_cellmath__32), .inst_cellmath__37__42__in1(inst_cellmath__28));
cynw_cm_float_mul_ieee_inst_cellmath__7_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I48 (.inst_cellmath__7_0_out0(inst_cellmath__7), .inst_cellmath__7_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__42_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I49 (.inst_cellmath__42_0_out0(inst_cellmath__42), .inst_cellmath__42_0_in0(inst_cellmath__7), .inst_cellmath__42_0_in1(inst_cellmath__6), .inst_cellmath__42_0_in2(inst_cellmath__5), .inst_cellmath__42_0_in3(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__52_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I50 (.inst_cellmath__52_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__52_0_in0(inst_cellmath__49), .inst_cellmath__52_0_in1({inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}), .inst_cellmath__52_0_in2(inst_cellmath__42), .inst_cellmath__52_0_in3({N470}), .inst_cellmath__52_0_in4({N469}));
cynw_cm_float_mul_ieee_inst_cellmath__47_0_bdw2876250654_bdw cynw_cm_float_mul_ieee_I51 (.inst_cellmath__47_0_out0(inst_cellmath__47), .inst_cellmath__47_0_in0(inst_cellmath__42), .inst_cellmath__47_0_in1(inst_cellmath__32), .inst_cellmath__47_0_in2(inst_cellmath__28), .inst_cellmath__47_0_in3(inst_cellmath__27), .inst_cellmath__47_0_in4(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__53_U_bdw2876250654_bdw cynw_cm_float_mul_ieee_I52 (.inst_cellmath__53_U_out0({x[22]}), .inst_cellmath__53_U_in0(inst_cellmath__49), .inst_cellmath__53_U_in1(inst_cellmath__47), .inst_cellmath__53_U_in2({inst_cellmath__45[22]}), .inst_cellmath__53_U_in3(inst_cellmath__44), .inst_cellmath__53_U_in4(inst_cellmath__26), .inst_cellmath__53_U_in5({inst_cellmath__25[46]}));
cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2876250654_bdw cynw_cm_float_mul_ieee_I53 (.inst_cellmath__53_M_out0({x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__53_M_in0(inst_cellmath__49), .inst_cellmath__53_M_in1(inst_cellmath__47), .inst_cellmath__53_M_in2({inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__53_M_in3(inst_cellmath__44), .inst_cellmath__53_M_in4(inst_cellmath__26), .inst_cellmath__53_M_in5({inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24]}), .inst_cellmath__53_M_in6(inst_cellmath__22), .inst_cellmath__53_M_in7(inst_cellmath__15), .inst_cellmath__53_M_in8({b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}), .inst_cellmath__53_M_in9({a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__17_0_bdw2876250654_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [7:0] inst_cellmath__17_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__17_0_I0 (.Y(N11), .A(inst_cellmath__17_0_in0[0]), .B(inst_cellmath__17_0_in0[1]));
NAND2XL inst_cellmath__17_0_I1 (.Y(N12), .A(inst_cellmath__17_0_in0[7]), .B(inst_cellmath__17_0_in0[6]));
NAND2XL inst_cellmath__17_0_I2 (.Y(N13), .A(inst_cellmath__17_0_in0[5]), .B(inst_cellmath__17_0_in0[4]));
NAND2XL inst_cellmath__17_0_I3 (.Y(N14), .A(inst_cellmath__17_0_in0[3]), .B(inst_cellmath__17_0_in0[2]));
NOR2XL inst_cellmath__17_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__17_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__17_0_I6 (.Y(inst_cellmath__17_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__19__2__bdw2876250654_bdw (
	inst_cellmath__19__2__out0,
	inst_cellmath__19__2__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__19__2__out0;
input [22:0] inst_cellmath__19__2__in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__19__2__I1 (.Y(N27), .A(inst_cellmath__19__2__in0[22]), .B(inst_cellmath__19__2__in0[21]));
NOR2XL inst_cellmath__19__2__I2 (.Y(N28), .A(inst_cellmath__19__2__in0[20]), .B(inst_cellmath__19__2__in0[19]));
NOR2XL inst_cellmath__19__2__I3 (.Y(N29), .A(inst_cellmath__19__2__in0[18]), .B(inst_cellmath__19__2__in0[17]));
NOR2XL inst_cellmath__19__2__I4 (.Y(N30), .A(inst_cellmath__19__2__in0[16]), .B(inst_cellmath__19__2__in0[15]));
NOR2XL inst_cellmath__19__2__I5 (.Y(N31), .A(inst_cellmath__19__2__in0[14]), .B(inst_cellmath__19__2__in0[13]));
NOR2XL inst_cellmath__19__2__I6 (.Y(N32), .A(inst_cellmath__19__2__in0[12]), .B(inst_cellmath__19__2__in0[11]));
NOR2XL inst_cellmath__19__2__I7 (.Y(N33), .A(inst_cellmath__19__2__in0[10]), .B(inst_cellmath__19__2__in0[9]));
NOR2XL inst_cellmath__19__2__I8 (.Y(N34), .A(inst_cellmath__19__2__in0[8]), .B(inst_cellmath__19__2__in0[7]));
NOR2XL inst_cellmath__19__2__I9 (.Y(N35), .A(inst_cellmath__19__2__in0[6]), .B(inst_cellmath__19__2__in0[5]));
NOR2XL inst_cellmath__19__2__I10 (.Y(N36), .A(inst_cellmath__19__2__in0[4]), .B(inst_cellmath__19__2__in0[3]));
NAND2XL inst_cellmath__19__2__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__19__2__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__19__2__I15 (.Y(N41), .A(N31), .B(N32));
NOR4XL inst_cellmath__19__2__I25 (.Y(N44), .A(inst_cellmath__19__2__in0[0]), .B(inst_cellmath__19__2__in0[1]), .C(inst_cellmath__19__2__in0[2]), .D(N39));
NOR2XL inst_cellmath__19__2__I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__19__2__I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__19__2__I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__19__2__I23 (.Y(inst_cellmath__19__2__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__21_0_bdw2876250654_bdw (
	inst_cellmath__21_0_out0,
	inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__21_0_out0;
input  inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1;
AND2XL inst_cellmath__21_0_I0 (.Y(inst_cellmath__21_0_out0), .A(inst_cellmath__21_0_in1), .B(inst_cellmath__21_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__13__1__bdw2876250654_bdw (
	inst_cellmath__13__1__out0,
	inst_cellmath__13__1__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__13__1__out0;
input [7:0] inst_cellmath__13__1__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2XL inst_cellmath__13__1__I0 (.Y(N11), .A(inst_cellmath__13__1__in0[0]), .B(inst_cellmath__13__1__in0[1]));
NOR2XL inst_cellmath__13__1__I1 (.Y(N12), .A(inst_cellmath__13__1__in0[7]), .B(inst_cellmath__13__1__in0[6]));
NOR2XL inst_cellmath__13__1__I2 (.Y(N13), .A(inst_cellmath__13__1__in0[5]), .B(inst_cellmath__13__1__in0[4]));
NOR2XL inst_cellmath__13__1__I3 (.Y(N14), .A(inst_cellmath__13__1__in0[3]), .B(inst_cellmath__13__1__in0[2]));
NAND2XL inst_cellmath__13__1__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__13__1__I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__13__1__I6 (.Y(inst_cellmath__13__1__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26__9__bdw2876250654_bdw (
	inst_cellmath__26__9__out0,
	inst_cellmath__26__9__in0,
	inst_cellmath__26__9__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__26__9__out0;
input  inst_cellmath__26__9__in0,
	inst_cellmath__26__9__in1;
AND2XL inst_cellmath__26__9__I0 (.Y(inst_cellmath__26__9__out0[0]), .A(inst_cellmath__26__9__in1), .B(inst_cellmath__26__9__in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__10_0_bdw2876250654_bdw (
	inst_cellmath__10_0_out0,
	inst_cellmath__10_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__10_0_out0;
input [7:0] inst_cellmath__10_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__10_0_I0 (.Y(N11), .A(inst_cellmath__10_0_in0[0]), .B(inst_cellmath__10_0_in0[1]));
NAND2XL inst_cellmath__10_0_I1 (.Y(N12), .A(inst_cellmath__10_0_in0[7]), .B(inst_cellmath__10_0_in0[6]));
NAND2XL inst_cellmath__10_0_I2 (.Y(N13), .A(inst_cellmath__10_0_in0[5]), .B(inst_cellmath__10_0_in0[4]));
NAND2XL inst_cellmath__10_0_I3 (.Y(N14), .A(inst_cellmath__10_0_in0[3]), .B(inst_cellmath__10_0_in0[2]));
NOR2XL inst_cellmath__10_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__10_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__10_0_I6 (.Y(inst_cellmath__10_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__12__0__bdw2876250654_bdw (
	inst_cellmath__12__0__out0,
	inst_cellmath__12__0__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__12__0__out0;
input [22:0] inst_cellmath__12__0__in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__12__0__I1 (.Y(N27), .A(inst_cellmath__12__0__in0[22]), .B(inst_cellmath__12__0__in0[21]));
NOR2XL inst_cellmath__12__0__I2 (.Y(N28), .A(inst_cellmath__12__0__in0[20]), .B(inst_cellmath__12__0__in0[19]));
NOR2XL inst_cellmath__12__0__I3 (.Y(N29), .A(inst_cellmath__12__0__in0[18]), .B(inst_cellmath__12__0__in0[17]));
NOR2XL inst_cellmath__12__0__I4 (.Y(N30), .A(inst_cellmath__12__0__in0[16]), .B(inst_cellmath__12__0__in0[15]));
NOR2XL inst_cellmath__12__0__I5 (.Y(N31), .A(inst_cellmath__12__0__in0[14]), .B(inst_cellmath__12__0__in0[13]));
NOR2XL inst_cellmath__12__0__I6 (.Y(N32), .A(inst_cellmath__12__0__in0[12]), .B(inst_cellmath__12__0__in0[11]));
NOR2XL inst_cellmath__12__0__I7 (.Y(N33), .A(inst_cellmath__12__0__in0[10]), .B(inst_cellmath__12__0__in0[9]));
NOR2XL inst_cellmath__12__0__I8 (.Y(N34), .A(inst_cellmath__12__0__in0[8]), .B(inst_cellmath__12__0__in0[7]));
NOR2XL inst_cellmath__12__0__I9 (.Y(N35), .A(inst_cellmath__12__0__in0[6]), .B(inst_cellmath__12__0__in0[5]));
NOR2XL inst_cellmath__12__0__I10 (.Y(N36), .A(inst_cellmath__12__0__in0[4]), .B(inst_cellmath__12__0__in0[3]));
NAND2XL inst_cellmath__12__0__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__12__0__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__12__0__I15 (.Y(N41), .A(N31), .B(N32));
NOR4X1 inst_cellmath__12__0__I25 (.Y(N44), .A(inst_cellmath__12__0__in0[0]), .B(inst_cellmath__12__0__in0[1]), .C(inst_cellmath__12__0__in0[2]), .D(N39));
NOR2XL inst_cellmath__12__0__I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__12__0__I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__12__0__I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__12__0__I23 (.Y(inst_cellmath__12__0__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__14_0_bdw2876250654_bdw (
	inst_cellmath__14_0_out0,
	inst_cellmath__14_0_in0,
	inst_cellmath__14_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__14_0_out0;
input  inst_cellmath__14_0_in0,
	inst_cellmath__14_0_in1;
AND2XL inst_cellmath__14_0_I0 (.Y(inst_cellmath__14_0_out0), .A(inst_cellmath__14_0_in1), .B(inst_cellmath__14_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__20__3__bdw2876250654_bdw (
	inst_cellmath__20__3__out0,
	inst_cellmath__20__3__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__20__3__out0;
input [7:0] inst_cellmath__20__3__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2XL inst_cellmath__20__3__I0 (.Y(N11), .A(inst_cellmath__20__3__in0[0]), .B(inst_cellmath__20__3__in0[1]));
NOR2XL inst_cellmath__20__3__I1 (.Y(N12), .A(inst_cellmath__20__3__in0[7]), .B(inst_cellmath__20__3__in0[6]));
NOR2XL inst_cellmath__20__3__I2 (.Y(N13), .A(inst_cellmath__20__3__in0[5]), .B(inst_cellmath__20__3__in0[4]));
NOR2XL inst_cellmath__20__3__I3 (.Y(N14), .A(inst_cellmath__20__3__in0[3]), .B(inst_cellmath__20__3__in0[2]));
NAND2XL inst_cellmath__20__3__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__20__3__I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__20__3__I6 (.Y(inst_cellmath__20__3__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26__8__bdw2876250654_bdw (
	inst_cellmath__26__8__out0,
	inst_cellmath__26__8__in0,
	inst_cellmath__26__8__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__26__8__out0;
input  inst_cellmath__26__8__in0,
	inst_cellmath__26__8__in1;
AND2XL inst_cellmath__26__8__I0 (.Y(inst_cellmath__26__8__out0[0]), .A(inst_cellmath__26__8__in0), .B(inst_cellmath__26__8__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__15_0_bdw2876250654_bdw (
	inst_cellmath__15_0_out0,
	inst_cellmath__15_0_in0,
	inst_cellmath__15_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__15_0_out0;
input  inst_cellmath__15_0_in0,
	inst_cellmath__15_0_in1;
NOR2BX1 inst_cellmath__15_0_I2 (.Y(inst_cellmath__15_0_out0), .AN(inst_cellmath__15_0_in1), .B(inst_cellmath__15_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__22_0_bdw2876250654_bdw (
	inst_cellmath__22_0_out0,
	inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__22_0_out0;
input  inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1;
NOR2BX1 inst_cellmath__22_0_I2 (.Y(inst_cellmath__22_0_out0), .AN(inst_cellmath__22_0_in1), .B(inst_cellmath__22_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26_1_bdw2876250654_bdw (
	inst_cellmath__26_1_out0,
	inst_cellmath__26_1_in0,
	inst_cellmath__26_1_in1,
	inst_cellmath__26_1_in2,
	inst_cellmath__26_1_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__26_1_out0;
input [0:0] inst_cellmath__26_1_in0,
	inst_cellmath__26_1_in1;
input  inst_cellmath__26_1_in2,
	inst_cellmath__26_1_in3;
OR4X1 inst_cellmath__26_1_I6 (.Y(inst_cellmath__26_1_out0), .A(inst_cellmath__26_1_in2), .B(inst_cellmath__26_1_in3), .C(inst_cellmath__26_1_in0[0]), .D(inst_cellmath__26_1_in1[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__23_0_bdw2876250654_bdw (
	inst_cellmath__23_0_out0,
	inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__23_0_out0;
input  inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1;
XOR2XL inst_cellmath__23_0_I0 (.Y(inst_cellmath__23_0_out0), .A(inst_cellmath__23_0_in1), .B(inst_cellmath__23_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__41_0_bdw2876250654_bdw (
	inst_cellmath__41_0_out0,
	inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2,
	inst_cellmath__41_0_in3,
	inst_cellmath__41_0_in4,
	inst_cellmath__41_0_in5
	); /* architecture "gate_level" */ 
output  inst_cellmath__41_0_out0;
input  inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2,
	inst_cellmath__41_0_in3,
	inst_cellmath__41_0_in4,
	inst_cellmath__41_0_in5;
wire N14,N16;
NAND2BXL inst_cellmath__41_0_I6 (.Y(N14), .AN(inst_cellmath__41_0_in4), .B(inst_cellmath__41_0_in2));
MX2XL inst_cellmath__41_0_I3 (.Y(N16), .A(N14), .B(inst_cellmath__41_0_in5), .S0(inst_cellmath__41_0_in3));
MX2XL inst_cellmath__41_0_I5 (.Y(inst_cellmath__41_0_out0), .A(inst_cellmath__41_0_in1), .B(N16), .S0(inst_cellmath__41_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__24_0_bdw2876250654_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1
	); /* architecture "gate_level" */ 
output [47:0] inst_cellmath__24_0_out0;
input [22:0] inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1;
wire N372,N381,N382,N384,N385,N386,N387 
	,N388,N389,N390,N391,N392,N393,N394,N395 
	,N396,N397,N398,N399,N400,N401,N402,N403 
	,N404,N405,N406,N407,N408,N409,N410,N411 
	,N412,N413,N414,N415,N416,N417,N418,N419 
	,N420,N421,N422,N423,N424,N425,N426,N427 
	,N428,N429,N438,N443,N444,N445,N446,N447 
	,N448,N449,N450,N451,N452,N453,N454,N455 
	,N456,N457,N458,N459,N460,N461,N462,N463 
	,N464,N465,N466,N467,N468,N469,N470,N471 
	,N472,N473,N474,N475,N476,N477,N478,N479 
	,N480,N481,N482,N483,N484,N485,N486,N487 
	,N488,N489,N490,N491,N492,N493,N502,N507 
	,N508,N509,N510,N511,N512,N513,N514,N515 
	,N516,N517,N518,N519,N520,N521,N522,N523 
	,N524,N525,N526,N527,N528,N529,N530,N531 
	,N532,N533,N534,N535,N536,N537,N538,N539 
	,N540,N541,N542,N543,N544,N545,N546,N547 
	,N548,N549,N550,N551,N552,N553,N554,N555 
	,N556,N557,N566,N567,N571,N572,N573,N574 
	,N575,N576,N577,N578,N579,N580,N581,N582 
	,N583,N584,N585,N586,N587,N588,N589,N590 
	,N591,N592,N593,N594,N595,N596,N597,N598 
	,N599,N600,N601,N602,N603,N604,N605,N606 
	,N607,N608,N609,N610,N611,N612,N613,N614 
	,N615,N616,N617,N618,N619,N620,N621,N630 
	,N631,N635,N636,N637,N638,N639,N640,N641 
	,N642,N643,N644,N645,N646,N647,N648,N649 
	,N650,N651,N652,N653,N654,N655,N656,N657 
	,N658,N659,N660,N661,N662,N663,N664,N665 
	,N666,N667,N668,N669,N670,N671,N672,N673 
	,N674,N675,N676,N677,N678,N679,N680,N681 
	,N682,N683,N684,N685,N694,N695,N699,N700 
	,N701,N702,N703,N704,N705,N706,N707,N708 
	,N709,N710,N711,N712,N713,N714,N715,N716 
	,N717,N718,N719,N720,N721,N722,N723,N724 
	,N725,N726,N727,N728,N729,N730,N731,N732 
	,N733,N734,N735,N736,N737,N738,N739,N740 
	,N741,N742,N743,N744,N745,N746,N747,N748 
	,N749,N758,N759,N763,N764,N765,N766,N767 
	,N768,N769,N770,N771,N772,N773,N774,N775 
	,N776,N777,N778,N779,N780,N781,N782,N783 
	,N784,N785,N786,N787,N788,N789,N790,N791 
	,N792,N793,N794,N795,N796,N797,N798,N799 
	,N800,N801,N802,N803,N804,N805,N806,N807 
	,N808,N809,N810,N811,N812,N813,N822,N823 
	,N827,N828,N829,N830,N831,N832,N833,N834 
	,N835,N836,N837,N838,N839,N840,N841,N842 
	,N843,N844,N845,N846,N847,N848,N849,N850 
	,N851,N852,N853,N854,N855,N856,N857,N858 
	,N859,N860,N861,N862,N863,N864,N865,N866 
	,N867,N868,N869,N870,N871,N872,N873,N874 
	,N875,N876,N877,N886,N887,N891,N892,N893 
	,N894,N895,N896,N897,N898,N899,N900,N901 
	,N902,N903,N904,N905,N906,N907,N908,N909 
	,N910,N911,N912,N913,N914,N915,N916,N917 
	,N918,N919,N920,N921,N922,N923,N924,N925 
	,N926,N927,N928,N929,N930,N931,N932,N933 
	,N934,N935,N936,N937,N938,N939,N940,N941 
	,N950,N955,N956,N957,N958,N959,N960,N961 
	,N962,N963,N964,N965,N966,N967,N968,N969 
	,N970,N971,N972,N973,N974,N975,N976,N977 
	,N978,N979,N980,N981,N982,N983,N984,N985 
	,N986,N987,N988,N989,N990,N991,N992,N993 
	,N994,N995,N996,N997,N998,N999,N1000,N1001 
	,N1002,N1003,N1004,N1005,N1014,N1019,N1020,N1021 
	,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029 
	,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037 
	,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045 
	,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053 
	,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061 
	,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069 
	,N1078,N1084,N1092,N1093,N1094,N1095,N1096,N1097 
	,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105 
	,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113 
	,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121 
	,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129 
	,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137 
	,N1138,N1140,N1144,N1212,N1213,N1214,N1215,N1216 
	,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224 
	,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232 
	,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240 
	,N1241,N1245,N1246,N1247,N1248,N1249,N1250,N1251 
	,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259 
	,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270 
	,N1271,N1275,N1276,N1277,N1278,N1279,N1280,N1281 
	,N1282,N1283,N1287,N1288,N1289,N1290,N1291,N1292 
	,N1293,N1294,N1295,N1296,N1297,N1301,N1302,N1303 
	,N1304,N1305,N1306,N1307,N1308,N1312,N1313,N1314 
	,N1315,N1319,N1320,N1321,N1322,N1323,N1324,N1325 
	,N1326,N1327,N1328,N1329,N1330,N1334,N1335,N1336 
	,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344 
	,N1345,N1349,N1350,N1351,N1352,N1353,N1354,N1355 
	,N1356,N1357,N1358,N1359,N1363,N1364,N1365,N1366 
	,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377 
	,N1378,N1379,N1380,N1384,N1385,N1386,N1387,N1391 
	,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399 
	,N1400,N1401,N1402,N1406,N1407,N1408,N1409,N1410 
	,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418 
	,N1419,N1420,N1424,N1425,N1426,N1427,N1428,N1429 
	,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437 
	,N1438,N1439,N1440,N1444,N1445,N1446,N1447,N1448 
	,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456 
	,N1457,N1458,N1459,N1460,N1464,N1465,N1466,N1467 
	,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478 
	,N1479,N1480,N1481,N1482,N1486,N1487,N1488,N1489 
	,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500 
	,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508 
	,N1509,N1510,N1514,N1515,N1516,N1517,N1521,N1522 
	,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530 
	,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538 
	,N1542,N1543,N1544,N1545,N1546,N1547,N1550,N1551 
	,N1552,N1553,N1554,N1555,N1559,N1560,N1561,N1562 
	,N1563,N1564,N1565,N1569,N1570,N1571,N1572,N1573 
	,N1574,N1577,N1578,N1579,N1580,N1581,N1582,N1583 
	,N1584,N1585,N1586,N1587,N1588,N1592,N1593,N1594 
	,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602 
	,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1613 
	,N1614,N1615,N1616,N1617,N1618,N1621,N1622,N1623 
	,N1624,N1625,N1626,N1627,N1628,N1632,N1633,N1634 
	,N1635,N1639,N1640,N1641,N1642,N1643,N1644,N1645 
	,N1646,N1647,N1648,N1649,N1650,N1651,N1655,N1656 
	,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1666 
	,N1667,N1668,N1672,N1673,N1674,N1675,N1679,N1680 
	,N1681,N1682,N1686,N1687,N1688,N1689,N1690,N1691 
	,N1692,N1693,N1694,N1695,N1696,N1697,N1701,N1702 
	,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1712 
	,N1713,N1714,N1715,N1716,N1720,N1721,N1722,N1723 
	,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734 
	,N1735,N1736,N1740,N1741,N1742,N1743,N1747,N1748 
	,N1749,N1750,N1751,N1752,N1755,N1756,N1757,N1761 
	,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769 
	,N1770,N1771,N1772,N1776,N1777,N1778,N1779,N1783 
	,N1784,N1785,N1786,N1787,N1788,N1791,N1792,N1796 
	,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804 
	,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812 
	,N1813,N1816,N1817,N1818,N1822,N1823,N1824,N1825 
	,N1826,N1827,N1828,N1829,N1830,N1834,N1835,N1836 
	,N1837,N1838,N1839,N1842,N1843,N1844,N1845,N1846 
	,N1847,N1848,N1849,N1853,N1854,N1855,N1856,N1857 
	,N1858,N1864,N1865,N1866,N1867,N1868,N1869,N1873 
	,N1874,N1875,N1876,N1877,N1878,N1881,N1882,N1886 
	,N1887,N1888,N1889,N1894,N1895,N1900,N1902,N1903 
	,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911 
	,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919 
	,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927 
	,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935 
	,N1936,N1937,N1940,N1950,N1958,N1970,N1982,N1998 
	,N2022,N2024,N2046,N2076,N2078,N2082,N2083,N2110 
	,N2148,N2150,N2154,N2155,N2202,N2204,N2218,N2221 
	,N2224,N2227,N2230,N2233,N2236,N2239,N2242,N2245 
	,N2248,N2251,N2254,N2257,N2260,N2263,N2266,N2287 
	,N2290,N2292,N2294,N2296,N2298,N2300,N2302,N2304 
	,N2306,N2308,N2310,N2312,N2314,N2316,N2318,N2320 
	,N2322,N2324,N2326,N2328,N2330,N2332,N2334,N2336 
	,N2338,N2340,N2342,N2344,N2346,N2349,N2355,N2363 
	,N2373,N2385,N2399,N2415,N2433,N2453,N2475,N2499 
	,N2525,N2553,N2583,N2615,N2649,N2685,N2723,N2763 
	,N2805,N2849,N2895,N2943,N2993,N3045,N3099,N3155 
	,N3213,N3737,N3964,N4191,N4418,N4645,N4872,N5099 
	,N5326,N5553,N5780,N6216,N6229,N6242,N6255,N6268 
	,N6281,N6294,N6307,N6320,N6333,N6346,N6359,N6372 
	,N6385,N6398,N6411,N6424,N6437,N6450,N6463,N6476 
	,N6489,N6502,N6515,N6528,N6541,N6554,N6567,N6580 
	,N6593,N6606,N6619,N6636,N6641,N6654,N6667,N6684 
	,N6689,N6702,N6715,N6728,N6741,N6754,N6767,N6780 
	,N6797,N6802,N6815,N6828,N6841,N6854,N6867,N6884 
	,N6889,N6902,N6915,N6928,N6945,N6950,N6963,N6976 
	,N6993,N6998,N7011,N7024,N7041,N7046,N7059,N7072 
	,N7085,N7102,N7107,N7120,N7137,N7142,N7155,N7172 
	,N7181,N7186,N7193,N7214,N7221,N7228,N7235,N7242 
	,N7249,N7256,N7263,N7270,N7277,N7284,N7291,N7298 
	,N7305,N7312,N7319,N7326,N7333,N7340,N7347,N7354 
	,N7361,N7368,N7375,N7670,N7671,N7672,N7673,N7674 
	,N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682 
	,N7683,N7684,N7685,N7686,N7687,N7688,N7689,N7690 
	,N7691,N7692,N7696,N7697,N7718,N7719,N7734,N7738 
	,N7740,N7741,N7763,N7785,N7807,N7829,N7841,N7863 
	,N7874,N7875,N7886,N7887,N7907,N7910,N7911,N7917 
	,N7918,N7928,N7929,N7940,N7949,N7950,N7964,N7965 
	,N7977,N7994,N7995,N8008,N8013,N8018,N8019,N8022 
	,N8028,N8035;
INVXL inst_cellmath__24_0_I3168 (.Y(N7670), .A(inst_cellmath__24_0_in1[0]));
INVXL inst_cellmath__24_0_I3169 (.Y(N7671), .A(inst_cellmath__24_0_in1[1]));
INVXL inst_cellmath__24_0_I3170 (.Y(N7672), .A(inst_cellmath__24_0_in1[2]));
INVXL inst_cellmath__24_0_I3171 (.Y(N7673), .A(inst_cellmath__24_0_in1[3]));
INVXL inst_cellmath__24_0_I3172 (.Y(N7674), .A(inst_cellmath__24_0_in1[4]));
INVXL inst_cellmath__24_0_I3173 (.Y(N7675), .A(inst_cellmath__24_0_in1[5]));
INVXL inst_cellmath__24_0_I3174 (.Y(N7676), .A(inst_cellmath__24_0_in1[6]));
INVXL inst_cellmath__24_0_I3175 (.Y(N7677), .A(inst_cellmath__24_0_in1[7]));
INVXL inst_cellmath__24_0_I3176 (.Y(N7678), .A(inst_cellmath__24_0_in1[8]));
INVXL inst_cellmath__24_0_I3177 (.Y(N7679), .A(inst_cellmath__24_0_in1[9]));
INVXL inst_cellmath__24_0_I3178 (.Y(N7680), .A(inst_cellmath__24_0_in1[10]));
INVXL inst_cellmath__24_0_I3179 (.Y(N7681), .A(inst_cellmath__24_0_in1[11]));
INVXL inst_cellmath__24_0_I3180 (.Y(N7682), .A(inst_cellmath__24_0_in1[12]));
INVXL inst_cellmath__24_0_I3181 (.Y(N7683), .A(inst_cellmath__24_0_in1[13]));
INVXL inst_cellmath__24_0_I3182 (.Y(N7684), .A(inst_cellmath__24_0_in1[14]));
INVXL inst_cellmath__24_0_I3183 (.Y(N7685), .A(inst_cellmath__24_0_in1[15]));
INVXL inst_cellmath__24_0_I3184 (.Y(N7686), .A(inst_cellmath__24_0_in1[16]));
INVXL inst_cellmath__24_0_I3185 (.Y(N7687), .A(inst_cellmath__24_0_in1[17]));
INVXL inst_cellmath__24_0_I3186 (.Y(N7688), .A(inst_cellmath__24_0_in1[18]));
INVXL inst_cellmath__24_0_I3187 (.Y(N7689), .A(inst_cellmath__24_0_in1[19]));
INVXL inst_cellmath__24_0_I3188 (.Y(N7690), .A(inst_cellmath__24_0_in1[20]));
INVXL inst_cellmath__24_0_I3189 (.Y(N7691), .A(inst_cellmath__24_0_in1[21]));
INVXL inst_cellmath__24_0_I3190 (.Y(N7692), .A(inst_cellmath__24_0_in1[22]));
INVXL inst_cellmath__24_0_I2222 (.Y(N372), .A(inst_cellmath__24_0_in0[0]));
NAND2X2 inst_cellmath__24_0_I3526 (.Y(N7696), .A(inst_cellmath__24_0_in0[1]), .B(N372));
INVX1 inst_cellmath__24_0_I3195 (.Y(N7697), .A(inst_cellmath__24_0_in0[1]));
XNOR2X1 addgen4_A_I2226 (.Y(N382), .A(N7670), .B(N7697));
OAI22XL addgen4_A_I2227 (.Y(N381), .A0(N382), .A1(N372), .B0(N7697), .B1(N7696));
XNOR2X1 addgen4_A_I2228 (.Y(N384), .A(N7671), .B(N7697));
OAI22XL addgen4_A_I2229 (.Y(N1903), .A0(N384), .A1(N372), .B0(N382), .B1(N7696));
XNOR2X1 addgen4_A_I2230 (.Y(N386), .A(N7672), .B(N7697));
OAI22XL addgen4_A_I2231 (.Y(N385), .A0(N386), .A1(N372), .B0(N384), .B1(N7696));
XNOR2X1 addgen4_A_I2232 (.Y(N388), .A(N7673), .B(N7697));
OAI22XL addgen4_A_I2233 (.Y(N387), .A0(N388), .A1(N372), .B0(N386), .B1(N7696));
XNOR2X1 addgen4_A_I2234 (.Y(N390), .A(N7674), .B(N7697));
OAI22XL addgen4_A_I2235 (.Y(N389), .A0(N390), .A1(N372), .B0(N388), .B1(N7696));
XNOR2X1 addgen4_A_I2236 (.Y(N392), .A(N7675), .B(N7697));
OAI22XL addgen4_A_I2237 (.Y(N391), .A0(N392), .A1(N372), .B0(N390), .B1(N7696));
XNOR2X1 addgen4_A_I2238 (.Y(N394), .A(N7676), .B(N7697));
OAI22XL addgen4_A_I2239 (.Y(N393), .A0(N394), .A1(N372), .B0(N392), .B1(N7696));
XNOR2X1 addgen4_A_I2240 (.Y(N396), .A(N7677), .B(N7697));
OAI22XL addgen4_A_I2241 (.Y(N395), .A0(N396), .A1(N372), .B0(N394), .B1(N7696));
XNOR2X1 addgen4_A_I2242 (.Y(N398), .A(N7678), .B(N7697));
OAI22XL addgen4_A_I2243 (.Y(N397), .A0(N398), .A1(N372), .B0(N396), .B1(N7696));
XNOR2X1 addgen4_A_I2244 (.Y(N400), .A(N7679), .B(N7697));
OAI22XL addgen4_A_I2245 (.Y(N399), .A0(N400), .A1(N372), .B0(N398), .B1(N7696));
XNOR2X1 addgen4_A_I2246 (.Y(N402), .A(N7680), .B(N7697));
OAI22XL addgen4_A_I2247 (.Y(N401), .A0(N402), .A1(N372), .B0(N400), .B1(N7696));
XNOR2X1 addgen4_A_I2248 (.Y(N404), .A(N7681), .B(N7697));
OAI22XL addgen4_A_I2249 (.Y(N403), .A0(N404), .A1(N372), .B0(N402), .B1(N7696));
XNOR2X1 addgen4_A_I2250 (.Y(N406), .A(N7682), .B(N7697));
OAI22XL addgen4_A_I2251 (.Y(N405), .A0(N406), .A1(N372), .B0(N404), .B1(N7696));
XNOR2X1 addgen4_A_I2252 (.Y(N408), .A(N7683), .B(N7697));
OAI22XL addgen4_A_I2253 (.Y(N407), .A0(N408), .A1(N372), .B0(N406), .B1(N7696));
XNOR2X1 addgen4_A_I2254 (.Y(N410), .A(N7684), .B(N7697));
OAI22XL addgen4_A_I2255 (.Y(N409), .A0(N410), .A1(N372), .B0(N408), .B1(N7696));
XNOR2X1 addgen4_A_I2256 (.Y(N412), .A(N7685), .B(N7697));
OAI22XL addgen4_A_I2257 (.Y(N411), .A0(N412), .A1(N372), .B0(N410), .B1(N7696));
XNOR2X1 addgen4_A_I2258 (.Y(N414), .A(N7686), .B(N7697));
OAI22XL addgen4_A_I2259 (.Y(N413), .A0(N414), .A1(N372), .B0(N412), .B1(N7696));
XNOR2X1 addgen4_A_I2260 (.Y(N416), .A(N7687), .B(N7697));
OAI22XL addgen4_A_I2261 (.Y(N415), .A0(N416), .A1(N372), .B0(N414), .B1(N7696));
XNOR2X1 addgen4_A_I2262 (.Y(N418), .A(N7688), .B(N7697));
OAI22XL addgen4_A_I2263 (.Y(N417), .A0(N418), .A1(N372), .B0(N416), .B1(N7696));
XNOR2X1 addgen4_A_I2264 (.Y(N420), .A(N7689), .B(N7697));
OAI22XL addgen4_A_I2265 (.Y(N419), .A0(N420), .A1(N372), .B0(N418), .B1(N7696));
XNOR2X1 addgen4_A_I2266 (.Y(N422), .A(N7690), .B(N7697));
OAI22XL addgen4_A_I2267 (.Y(N421), .A0(N422), .A1(N372), .B0(N420), .B1(N7696));
XNOR2X1 addgen4_A_I2268 (.Y(N424), .A(N7691), .B(N7697));
OAI22XL addgen4_A_I2269 (.Y(N423), .A0(N424), .A1(N372), .B0(N422), .B1(N7696));
XNOR2X1 addgen4_A_I2270 (.Y(N426), .A(N7692), .B(N7697));
OAI22XL addgen4_A_I2271 (.Y(N425), .A0(N426), .A1(N372), .B0(N424), .B1(N7696));
INVXL addgen4_A_I2272 (.Y(N428), .A(N7697));
OAI22XL addgen4_A_I2273 (.Y(N427), .A0(N428), .A1(N372), .B0(N426), .B1(N7696));
MXI2XL inst_cellmath__24_0_I113 (.Y(N429), .A(N7696), .B(N372), .S0(N428));
XNOR2X1 enc3_A_I2274 (.Y(N438), .A(inst_cellmath__24_0_in0[2]), .B(inst_cellmath__24_0_in0[1]));
XOR2XL enc3_A_I2275 (.Y(N3737), .A(inst_cellmath__24_0_in0[3]), .B(inst_cellmath__24_0_in0[1]));
NAND2X2 inst_cellmath__24_0_I3568 (.Y(N7718), .A(N3737), .B(N438));
INVX1 inst_cellmath__24_0_I3217 (.Y(N7719), .A(inst_cellmath__24_0_in0[3]));
NAND2XL inst_cellmath__24_0_I119 (.Y(N443), .A(inst_cellmath__24_0_in0[1]), .B(inst_cellmath__24_0_in0[2]));
AND2XL inst_cellmath__24_0_I120 (.Y(N444), .A(inst_cellmath__24_0_in0[3]), .B(N443));
XNOR2X1 addgen4_A_I2278 (.Y(N446), .A(N7670), .B(N7719));
OAI22XL addgen4_A_I2279 (.Y(N445), .A0(N446), .A1(N438), .B0(N7719), .B1(N7718));
XNOR2X1 addgen4_A_I2280 (.Y(N448), .A(N7671), .B(N7719));
OAI22XL addgen4_A_I2281 (.Y(N447), .A0(N448), .A1(N438), .B0(N446), .B1(N7718));
XNOR2X1 addgen4_A_I2282 (.Y(N450), .A(N7672), .B(N7719));
OAI22XL addgen4_A_I2283 (.Y(N449), .A0(N450), .A1(N438), .B0(N448), .B1(N7718));
XNOR2X1 addgen4_A_I2284 (.Y(N452), .A(N7673), .B(N7719));
OAI22XL addgen4_A_I2285 (.Y(N451), .A0(N452), .A1(N438), .B0(N450), .B1(N7718));
XNOR2X1 addgen4_A_I2286 (.Y(N454), .A(N7674), .B(N7719));
OAI22XL addgen4_A_I2287 (.Y(N453), .A0(N454), .A1(N438), .B0(N452), .B1(N7718));
XNOR2X1 addgen4_A_I2288 (.Y(N456), .A(N7675), .B(N7719));
OAI22XL addgen4_A_I2289 (.Y(N455), .A0(N456), .A1(N438), .B0(N454), .B1(N7718));
XNOR2X1 addgen4_A_I2290 (.Y(N458), .A(N7676), .B(N7719));
OAI22XL addgen4_A_I2291 (.Y(N457), .A0(N458), .A1(N438), .B0(N456), .B1(N7718));
XNOR2X1 addgen4_A_I2292 (.Y(N460), .A(N7677), .B(N7719));
OAI22XL addgen4_A_I2293 (.Y(N459), .A0(N460), .A1(N438), .B0(N458), .B1(N7718));
XNOR2X1 addgen4_A_I2294 (.Y(N462), .A(N7678), .B(N7719));
OAI22XL addgen4_A_I2295 (.Y(N461), .A0(N462), .A1(N438), .B0(N460), .B1(N7718));
XNOR2X1 addgen4_A_I2296 (.Y(N464), .A(N7679), .B(N7719));
OAI22XL addgen4_A_I2297 (.Y(N463), .A0(N464), .A1(N438), .B0(N462), .B1(N7718));
XNOR2X1 addgen4_A_I2298 (.Y(N466), .A(N7680), .B(N7719));
OAI22XL addgen4_A_I2299 (.Y(N465), .A0(N466), .A1(N438), .B0(N464), .B1(N7718));
XNOR2X1 addgen4_A_I2300 (.Y(N468), .A(N7681), .B(N7719));
OAI22XL addgen4_A_I2301 (.Y(N467), .A0(N468), .A1(N438), .B0(N466), .B1(N7718));
XNOR2X1 addgen4_A_I2302 (.Y(N470), .A(N7682), .B(N7719));
OAI22XL addgen4_A_I2303 (.Y(N469), .A0(N470), .A1(N438), .B0(N468), .B1(N7718));
XNOR2X1 addgen4_A_I2304 (.Y(N472), .A(N7683), .B(N7719));
OAI22XL addgen4_A_I2305 (.Y(N471), .A0(N472), .A1(N438), .B0(N470), .B1(N7718));
XNOR2X1 addgen4_A_I2306 (.Y(N474), .A(N7684), .B(N7719));
OAI22XL addgen4_A_I2307 (.Y(N473), .A0(N474), .A1(N438), .B0(N472), .B1(N7718));
XNOR2X1 addgen4_A_I2308 (.Y(N476), .A(N7685), .B(N7719));
OAI22XL addgen4_A_I2309 (.Y(N475), .A0(N476), .A1(N438), .B0(N474), .B1(N7718));
XNOR2X1 addgen4_A_I2310 (.Y(N478), .A(N7686), .B(N7719));
OAI22XL addgen4_A_I2311 (.Y(N477), .A0(N478), .A1(N438), .B0(N476), .B1(N7718));
XNOR2X1 addgen4_A_I2312 (.Y(N480), .A(N7687), .B(N7719));
OAI22XL addgen4_A_I2313 (.Y(N479), .A0(N480), .A1(N438), .B0(N478), .B1(N7718));
XNOR2X1 addgen4_A_I2314 (.Y(N482), .A(N7688), .B(N7719));
OAI22XL addgen4_A_I2315 (.Y(N481), .A0(N482), .A1(N438), .B0(N480), .B1(N7718));
XNOR2X1 addgen4_A_I2316 (.Y(N484), .A(N7689), .B(N7719));
OAI22XL addgen4_A_I2317 (.Y(N483), .A0(N484), .A1(N438), .B0(N482), .B1(N7718));
XNOR2X1 addgen4_A_I2318 (.Y(N486), .A(N7690), .B(N7719));
OAI22XL addgen4_A_I2319 (.Y(N485), .A0(N486), .A1(N438), .B0(N484), .B1(N7718));
XNOR2X1 addgen4_A_I2320 (.Y(N488), .A(N7691), .B(N7719));
OAI22XL addgen4_A_I2321 (.Y(N487), .A0(N488), .A1(N438), .B0(N486), .B1(N7718));
XNOR2X1 addgen4_A_I2322 (.Y(N490), .A(N7692), .B(N7719));
OAI22XL addgen4_A_I2323 (.Y(N489), .A0(N490), .A1(N438), .B0(N488), .B1(N7718));
INVXL addgen4_A_I2324 (.Y(N492), .A(N7719));
OAI22XL addgen4_A_I2325 (.Y(N491), .A0(N492), .A1(N438), .B0(N490), .B1(N7718));
MXI2XL inst_cellmath__24_0_I145 (.Y(N493), .A(N7718), .B(N438), .S0(N492));
XNOR2X1 enc3_A_I2326 (.Y(N502), .A(inst_cellmath__24_0_in0[4]), .B(inst_cellmath__24_0_in0[3]));
XOR2XL enc3_A_I2327 (.Y(N3964), .A(inst_cellmath__24_0_in0[5]), .B(inst_cellmath__24_0_in0[3]));
AND2XL inst_cellmath__24_0_I3529 (.Y(N7734), .A(N3964), .B(N502));
INVXL inst_cellmath__24_0_I3238 (.Y(N7740), .A(N7734));
INVXL inst_cellmath__24_0_I3236 (.Y(N7738), .A(N7734));
INVX1 inst_cellmath__24_0_I3239 (.Y(N7741), .A(inst_cellmath__24_0_in0[5]));
NAND2XL inst_cellmath__24_0_I151 (.Y(N507), .A(inst_cellmath__24_0_in0[3]), .B(inst_cellmath__24_0_in0[4]));
AND2XL inst_cellmath__24_0_I152 (.Y(N508), .A(inst_cellmath__24_0_in0[5]), .B(N507));
XNOR2X1 addgen4_A_I2330 (.Y(N510), .A(N7670), .B(N7741));
OAI22XL addgen4_A_I2331 (.Y(N509), .A0(N510), .A1(N502), .B0(N7741), .B1(N7740));
XNOR2X1 addgen4_A_I2332 (.Y(N512), .A(N7671), .B(N7741));
OAI22XL addgen4_A_I2333 (.Y(N511), .A0(N512), .A1(N502), .B0(N510), .B1(N7740));
XNOR2X1 addgen4_A_I2334 (.Y(N514), .A(N7672), .B(N7741));
OAI22XL addgen4_A_I2335 (.Y(N513), .A0(N514), .A1(N502), .B0(N512), .B1(N7740));
XNOR2X1 addgen4_A_I2336 (.Y(N516), .A(N7673), .B(N7741));
OAI22XL addgen4_A_I2337 (.Y(N515), .A0(N516), .A1(N502), .B0(N514), .B1(N7740));
XNOR2X1 addgen4_A_I2338 (.Y(N518), .A(N7674), .B(N7741));
OAI22XL addgen4_A_I2339 (.Y(N517), .A0(N518), .A1(N502), .B0(N516), .B1(N7740));
XNOR2X1 addgen4_A_I2340 (.Y(N520), .A(N7675), .B(N7741));
OAI22XL addgen4_A_I2341 (.Y(N519), .A0(N520), .A1(N502), .B0(N518), .B1(N7738));
XNOR2X1 addgen4_A_I2342 (.Y(N522), .A(N7676), .B(N7741));
OAI22XL addgen4_A_I2343 (.Y(N521), .A0(N522), .A1(N502), .B0(N520), .B1(N7738));
XNOR2X1 addgen4_A_I2344 (.Y(N524), .A(N7677), .B(N7741));
OAI22XL addgen4_A_I2345 (.Y(N523), .A0(N524), .A1(N502), .B0(N522), .B1(N7738));
XNOR2X1 addgen4_A_I2346 (.Y(N526), .A(N7678), .B(N7741));
OAI22XL addgen4_A_I2347 (.Y(N525), .A0(N526), .A1(N502), .B0(N524), .B1(N7738));
XNOR2X1 addgen4_A_I2348 (.Y(N528), .A(N7679), .B(N7741));
OAI22XL addgen4_A_I2349 (.Y(N527), .A0(N528), .A1(N502), .B0(N526), .B1(N7738));
XNOR2X1 addgen4_A_I2350 (.Y(N530), .A(N7680), .B(N7741));
OAI22XL addgen4_A_I2351 (.Y(N529), .A0(N530), .A1(N502), .B0(N528), .B1(N7738));
XNOR2X1 addgen4_A_I2352 (.Y(N532), .A(N7681), .B(N7741));
OAI22XL addgen4_A_I2353 (.Y(N531), .A0(N532), .A1(N502), .B0(N530), .B1(N7738));
XNOR2X1 addgen4_A_I2354 (.Y(N534), .A(N7682), .B(N7741));
OAI22XL addgen4_A_I2355 (.Y(N533), .A0(N534), .A1(N502), .B0(N532), .B1(N7738));
XNOR2X1 addgen4_A_I2356 (.Y(N536), .A(N7683), .B(N7741));
OAI22XL addgen4_A_I2357 (.Y(N535), .A0(N536), .A1(N502), .B0(N534), .B1(N7738));
XNOR2X1 addgen4_A_I2358 (.Y(N538), .A(N7684), .B(N7741));
OAI22XL addgen4_A_I2359 (.Y(N537), .A0(N538), .A1(N502), .B0(N536), .B1(N7738));
XNOR2X1 addgen4_A_I2360 (.Y(N540), .A(N7685), .B(N7741));
OAI22XL addgen4_A_I2361 (.Y(N539), .A0(N540), .A1(N502), .B0(N538), .B1(N7740));
XNOR2X1 addgen4_A_I2362 (.Y(N542), .A(N7686), .B(N7741));
OAI22XL addgen4_A_I2363 (.Y(N541), .A0(N542), .A1(N502), .B0(N540), .B1(N7740));
XNOR2X1 addgen4_A_I2364 (.Y(N544), .A(N7687), .B(N7741));
OAI22XL addgen4_A_I2365 (.Y(N543), .A0(N544), .A1(N502), .B0(N542), .B1(N7740));
XNOR2X1 addgen4_A_I2366 (.Y(N546), .A(N7688), .B(N7741));
OAI22XL addgen4_A_I2367 (.Y(N545), .A0(N546), .A1(N502), .B0(N544), .B1(N7740));
XNOR2X1 addgen4_A_I2368 (.Y(N548), .A(N7689), .B(N7741));
OAI22XL addgen4_A_I2369 (.Y(N547), .A0(N548), .A1(N502), .B0(N546), .B1(N7740));
XNOR2X1 addgen4_A_I2370 (.Y(N550), .A(N7690), .B(N7741));
OAI22XL addgen4_A_I2371 (.Y(N549), .A0(N550), .A1(N502), .B0(N548), .B1(N7740));
XNOR2X1 addgen4_A_I2372 (.Y(N552), .A(N7691), .B(N7741));
OAI22XL addgen4_A_I2373 (.Y(N551), .A0(N552), .A1(N502), .B0(N550), .B1(N7740));
XNOR2X1 addgen4_A_I2374 (.Y(N554), .A(N7692), .B(N7741));
OAI22XL addgen4_A_I2375 (.Y(N553), .A0(N554), .A1(N502), .B0(N552), .B1(N7740));
INVXL addgen4_A_I2376 (.Y(N556), .A(N7741));
OAI22XL addgen4_A_I2377 (.Y(N555), .A0(N556), .A1(N502), .B0(N554), .B1(N7740));
MXI2XL inst_cellmath__24_0_I177 (.Y(N557), .A(N7740), .B(N502), .S0(N556));
XNOR2X1 enc3_A_I2378 (.Y(N566), .A(inst_cellmath__24_0_in0[6]), .B(inst_cellmath__24_0_in0[5]));
XOR2XL enc3_A_I2379 (.Y(N4191), .A(inst_cellmath__24_0_in0[7]), .B(inst_cellmath__24_0_in0[5]));
NAND2X2 enc3_A_I2381 (.Y(N567), .A(N4191), .B(N566));
INVX1 inst_cellmath__24_0_I3261 (.Y(N7763), .A(inst_cellmath__24_0_in0[7]));
NAND2XL inst_cellmath__24_0_I183 (.Y(N571), .A(inst_cellmath__24_0_in0[5]), .B(inst_cellmath__24_0_in0[6]));
AND2XL inst_cellmath__24_0_I184 (.Y(N572), .A(inst_cellmath__24_0_in0[7]), .B(N571));
XNOR2X1 addgen4_A_I2382 (.Y(N574), .A(N7670), .B(N7763));
OAI22XL addgen4_A_I2383 (.Y(N573), .A0(N574), .A1(N566), .B0(N7763), .B1(N567));
XNOR2X1 addgen4_A_I2384 (.Y(N576), .A(N7671), .B(N7763));
OAI22XL addgen4_A_I2385 (.Y(N575), .A0(N576), .A1(N566), .B0(N574), .B1(N567));
XNOR2X1 addgen4_A_I2386 (.Y(N578), .A(N7672), .B(N7763));
OAI22XL addgen4_A_I2387 (.Y(N577), .A0(N578), .A1(N566), .B0(N576), .B1(N567));
XNOR2X1 addgen4_A_I2388 (.Y(N580), .A(N7673), .B(N7763));
OAI22XL addgen4_A_I2389 (.Y(N579), .A0(N580), .A1(N566), .B0(N578), .B1(N567));
XNOR2X1 addgen4_A_I2390 (.Y(N582), .A(N7674), .B(N7763));
OAI22XL addgen4_A_I2391 (.Y(N581), .A0(N582), .A1(N566), .B0(N580), .B1(N567));
XNOR2X1 addgen4_A_I2392 (.Y(N584), .A(N7675), .B(N7763));
OAI22XL addgen4_A_I2393 (.Y(N583), .A0(N584), .A1(N566), .B0(N582), .B1(N567));
XNOR2X1 addgen4_A_I2394 (.Y(N586), .A(N7676), .B(N7763));
OAI22XL addgen4_A_I2395 (.Y(N585), .A0(N586), .A1(N566), .B0(N584), .B1(N567));
XNOR2X1 addgen4_A_I2396 (.Y(N588), .A(N7677), .B(N7763));
OAI22XL addgen4_A_I2397 (.Y(N587), .A0(N588), .A1(N566), .B0(N586), .B1(N567));
XNOR2X1 addgen4_A_I2398 (.Y(N590), .A(N7678), .B(N7763));
OAI22XL addgen4_A_I2399 (.Y(N589), .A0(N590), .A1(N566), .B0(N588), .B1(N567));
XNOR2X1 addgen4_A_I2400 (.Y(N592), .A(N7679), .B(N7763));
OAI22XL addgen4_A_I2401 (.Y(N591), .A0(N592), .A1(N566), .B0(N590), .B1(N567));
XNOR2X1 addgen4_A_I2402 (.Y(N594), .A(N7680), .B(N7763));
OAI22XL addgen4_A_I2403 (.Y(N593), .A0(N594), .A1(N566), .B0(N592), .B1(N567));
XNOR2X1 addgen4_A_I2404 (.Y(N596), .A(N7681), .B(N7763));
OAI22XL addgen4_A_I2405 (.Y(N595), .A0(N596), .A1(N566), .B0(N594), .B1(N567));
XNOR2X1 addgen4_A_I2406 (.Y(N598), .A(N7682), .B(N7763));
OAI22XL addgen4_A_I2407 (.Y(N597), .A0(N598), .A1(N566), .B0(N596), .B1(N567));
XNOR2X1 addgen4_A_I2408 (.Y(N600), .A(N7683), .B(N7763));
OAI22XL addgen4_A_I2409 (.Y(N599), .A0(N600), .A1(N566), .B0(N598), .B1(N567));
XNOR2X1 addgen4_A_I2410 (.Y(N602), .A(N7684), .B(N7763));
OAI22XL addgen4_A_I2411 (.Y(N601), .A0(N602), .A1(N566), .B0(N600), .B1(N567));
XNOR2X1 addgen4_A_I2412 (.Y(N604), .A(N7685), .B(N7763));
OAI22XL addgen4_A_I2413 (.Y(N603), .A0(N604), .A1(N566), .B0(N602), .B1(N567));
XNOR2X1 addgen4_A_I2414 (.Y(N606), .A(N7686), .B(N7763));
OAI22XL addgen4_A_I2415 (.Y(N605), .A0(N606), .A1(N566), .B0(N604), .B1(N567));
XNOR2X1 addgen4_A_I2416 (.Y(N608), .A(N7687), .B(N7763));
OAI22XL addgen4_A_I2417 (.Y(N607), .A0(N608), .A1(N566), .B0(N606), .B1(N567));
XNOR2X1 addgen4_A_I2418 (.Y(N610), .A(N7688), .B(N7763));
OAI22XL addgen4_A_I2419 (.Y(N609), .A0(N610), .A1(N566), .B0(N608), .B1(N567));
XNOR2X1 addgen4_A_I2420 (.Y(N612), .A(N7689), .B(N7763));
OAI22XL addgen4_A_I2421 (.Y(N611), .A0(N612), .A1(N566), .B0(N610), .B1(N567));
XNOR2X1 addgen4_A_I2422 (.Y(N614), .A(N7690), .B(N7763));
OAI22XL addgen4_A_I2423 (.Y(N613), .A0(N614), .A1(N566), .B0(N612), .B1(N567));
XNOR2X1 addgen4_A_I2424 (.Y(N616), .A(N7691), .B(N7763));
OAI22XL addgen4_A_I2425 (.Y(N615), .A0(N616), .A1(N566), .B0(N614), .B1(N567));
XNOR2X1 addgen4_A_I2426 (.Y(N618), .A(N7692), .B(N7763));
OAI22XL addgen4_A_I2427 (.Y(N617), .A0(N618), .A1(N566), .B0(N616), .B1(N567));
INVXL addgen4_A_I2428 (.Y(N620), .A(N7763));
OAI22XL addgen4_A_I2429 (.Y(N619), .A0(N620), .A1(N566), .B0(N618), .B1(N567));
MXI2XL inst_cellmath__24_0_I209 (.Y(N621), .A(N567), .B(N566), .S0(N620));
XNOR2X1 enc3_A_I2430 (.Y(N630), .A(inst_cellmath__24_0_in0[8]), .B(inst_cellmath__24_0_in0[7]));
XOR2XL enc3_A_I2431 (.Y(N4418), .A(inst_cellmath__24_0_in0[9]), .B(inst_cellmath__24_0_in0[7]));
NAND2X2 enc3_A_I2433 (.Y(N631), .A(N4418), .B(N630));
INVX1 inst_cellmath__24_0_I3283 (.Y(N7785), .A(inst_cellmath__24_0_in0[9]));
NAND2XL inst_cellmath__24_0_I215 (.Y(N635), .A(inst_cellmath__24_0_in0[7]), .B(inst_cellmath__24_0_in0[8]));
AND2XL inst_cellmath__24_0_I216 (.Y(N636), .A(inst_cellmath__24_0_in0[9]), .B(N635));
XNOR2X1 addgen4_A_I2434 (.Y(N638), .A(N7670), .B(N7785));
OAI22XL addgen4_A_I2435 (.Y(N637), .A0(N638), .A1(N630), .B0(N7785), .B1(N631));
XNOR2X1 addgen4_A_I2436 (.Y(N640), .A(N7671), .B(N7785));
OAI22XL addgen4_A_I2437 (.Y(N639), .A0(N640), .A1(N630), .B0(N638), .B1(N631));
XNOR2X1 addgen4_A_I2438 (.Y(N642), .A(N7672), .B(N7785));
OAI22XL addgen4_A_I2439 (.Y(N641), .A0(N642), .A1(N630), .B0(N640), .B1(N631));
XNOR2X1 addgen4_A_I2440 (.Y(N644), .A(N7673), .B(N7785));
OAI22XL addgen4_A_I2441 (.Y(N643), .A0(N644), .A1(N630), .B0(N642), .B1(N631));
XNOR2X1 addgen4_A_I2442 (.Y(N646), .A(N7674), .B(N7785));
OAI22XL addgen4_A_I2443 (.Y(N645), .A0(N646), .A1(N630), .B0(N644), .B1(N631));
XNOR2X1 addgen4_A_I2444 (.Y(N648), .A(N7675), .B(N7785));
OAI22XL addgen4_A_I2445 (.Y(N647), .A0(N648), .A1(N630), .B0(N646), .B1(N631));
XNOR2X1 addgen4_A_I2446 (.Y(N650), .A(N7676), .B(N7785));
OAI22XL addgen4_A_I2447 (.Y(N649), .A0(N650), .A1(N630), .B0(N648), .B1(N631));
XNOR2X1 addgen4_A_I2448 (.Y(N652), .A(N7677), .B(N7785));
OAI22XL addgen4_A_I2449 (.Y(N651), .A0(N652), .A1(N630), .B0(N650), .B1(N631));
XNOR2X1 addgen4_A_I2450 (.Y(N654), .A(N7678), .B(N7785));
OAI22XL addgen4_A_I2451 (.Y(N653), .A0(N654), .A1(N630), .B0(N652), .B1(N631));
XNOR2X1 addgen4_A_I2452 (.Y(N656), .A(N7679), .B(N7785));
OAI22XL addgen4_A_I2453 (.Y(N655), .A0(N656), .A1(N630), .B0(N654), .B1(N631));
XNOR2X1 addgen4_A_I2454 (.Y(N658), .A(N7680), .B(N7785));
OAI22XL addgen4_A_I2455 (.Y(N657), .A0(N658), .A1(N630), .B0(N656), .B1(N631));
XNOR2X1 addgen4_A_I2456 (.Y(N660), .A(N7681), .B(N7785));
OAI22XL addgen4_A_I2457 (.Y(N659), .A0(N660), .A1(N630), .B0(N658), .B1(N631));
XNOR2X1 addgen4_A_I2458 (.Y(N662), .A(N7682), .B(N7785));
OAI22XL addgen4_A_I2459 (.Y(N661), .A0(N662), .A1(N630), .B0(N660), .B1(N631));
XNOR2X1 addgen4_A_I2460 (.Y(N664), .A(N7683), .B(N7785));
OAI22XL addgen4_A_I2461 (.Y(N663), .A0(N664), .A1(N630), .B0(N662), .B1(N631));
XNOR2X1 addgen4_A_I2462 (.Y(N666), .A(N7684), .B(N7785));
OAI22XL addgen4_A_I2463 (.Y(N665), .A0(N666), .A1(N630), .B0(N664), .B1(N631));
XNOR2X1 addgen4_A_I2464 (.Y(N668), .A(N7685), .B(N7785));
OAI22XL addgen4_A_I2465 (.Y(N667), .A0(N668), .A1(N630), .B0(N666), .B1(N631));
XNOR2X1 addgen4_A_I2466 (.Y(N670), .A(N7686), .B(N7785));
OAI22XL addgen4_A_I2467 (.Y(N669), .A0(N670), .A1(N630), .B0(N668), .B1(N631));
XNOR2X1 addgen4_A_I2468 (.Y(N672), .A(N7687), .B(N7785));
OAI22XL addgen4_A_I2469 (.Y(N671), .A0(N672), .A1(N630), .B0(N670), .B1(N631));
XNOR2X1 addgen4_A_I2470 (.Y(N674), .A(N7688), .B(N7785));
OAI22XL addgen4_A_I2471 (.Y(N673), .A0(N674), .A1(N630), .B0(N672), .B1(N631));
XNOR2X1 addgen4_A_I2472 (.Y(N676), .A(N7689), .B(N7785));
OAI22XL addgen4_A_I2473 (.Y(N675), .A0(N676), .A1(N630), .B0(N674), .B1(N631));
XNOR2X1 addgen4_A_I2474 (.Y(N678), .A(N7690), .B(N7785));
OAI22XL addgen4_A_I2475 (.Y(N677), .A0(N678), .A1(N630), .B0(N676), .B1(N631));
XNOR2X1 addgen4_A_I2476 (.Y(N680), .A(N7691), .B(N7785));
OAI22XL addgen4_A_I2477 (.Y(N679), .A0(N680), .A1(N630), .B0(N678), .B1(N631));
XNOR2X1 addgen4_A_I2478 (.Y(N682), .A(N7692), .B(N7785));
OAI22XL addgen4_A_I2479 (.Y(N681), .A0(N682), .A1(N630), .B0(N680), .B1(N631));
INVXL addgen4_A_I2480 (.Y(N684), .A(N7785));
OAI22XL addgen4_A_I2481 (.Y(N683), .A0(N684), .A1(N630), .B0(N682), .B1(N631));
MXI2XL inst_cellmath__24_0_I241 (.Y(N685), .A(N631), .B(N630), .S0(N684));
XNOR2X1 enc3_A_I2482 (.Y(N694), .A(inst_cellmath__24_0_in0[10]), .B(inst_cellmath__24_0_in0[9]));
XOR2XL enc3_A_I2483 (.Y(N4645), .A(inst_cellmath__24_0_in0[11]), .B(inst_cellmath__24_0_in0[9]));
NAND2X2 enc3_A_I2485 (.Y(N695), .A(N4645), .B(N694));
INVX1 inst_cellmath__24_0_I3305 (.Y(N7807), .A(inst_cellmath__24_0_in0[11]));
NAND2XL inst_cellmath__24_0_I247 (.Y(N699), .A(inst_cellmath__24_0_in0[9]), .B(inst_cellmath__24_0_in0[10]));
AND2XL inst_cellmath__24_0_I248 (.Y(N700), .A(inst_cellmath__24_0_in0[11]), .B(N699));
XNOR2X1 addgen4_A_I2486 (.Y(N702), .A(N7670), .B(N7807));
OAI22XL addgen4_A_I2487 (.Y(N701), .A0(N702), .A1(N694), .B0(N7807), .B1(N695));
XNOR2X1 addgen4_A_I2488 (.Y(N704), .A(N7671), .B(N7807));
OAI22XL addgen4_A_I2489 (.Y(N703), .A0(N704), .A1(N694), .B0(N702), .B1(N695));
XNOR2X1 addgen4_A_I2490 (.Y(N706), .A(N7672), .B(N7807));
OAI22XL addgen4_A_I2491 (.Y(N705), .A0(N706), .A1(N694), .B0(N704), .B1(N695));
XNOR2X1 addgen4_A_I2492 (.Y(N708), .A(N7673), .B(N7807));
OAI22XL addgen4_A_I2493 (.Y(N707), .A0(N708), .A1(N694), .B0(N706), .B1(N695));
XNOR2X1 addgen4_A_I2494 (.Y(N710), .A(N7674), .B(N7807));
OAI22XL addgen4_A_I2495 (.Y(N709), .A0(N710), .A1(N694), .B0(N708), .B1(N695));
XNOR2X1 addgen4_A_I2496 (.Y(N712), .A(N7675), .B(N7807));
OAI22XL addgen4_A_I2497 (.Y(N711), .A0(N712), .A1(N694), .B0(N710), .B1(N695));
XNOR2X1 addgen4_A_I2498 (.Y(N714), .A(N7676), .B(N7807));
OAI22XL addgen4_A_I2499 (.Y(N713), .A0(N714), .A1(N694), .B0(N712), .B1(N695));
XNOR2X1 addgen4_A_I2500 (.Y(N716), .A(N7677), .B(N7807));
OAI22XL addgen4_A_I2501 (.Y(N715), .A0(N716), .A1(N694), .B0(N714), .B1(N695));
XNOR2X1 addgen4_A_I2502 (.Y(N718), .A(N7678), .B(N7807));
OAI22XL addgen4_A_I2503 (.Y(N717), .A0(N718), .A1(N694), .B0(N716), .B1(N695));
XNOR2X1 addgen4_A_I2504 (.Y(N720), .A(N7679), .B(N7807));
OAI22XL addgen4_A_I2505 (.Y(N719), .A0(N720), .A1(N694), .B0(N718), .B1(N695));
XNOR2X1 addgen4_A_I2506 (.Y(N722), .A(N7680), .B(N7807));
OAI22XL addgen4_A_I2507 (.Y(N721), .A0(N722), .A1(N694), .B0(N720), .B1(N695));
XNOR2X1 addgen4_A_I2508 (.Y(N724), .A(N7681), .B(N7807));
OAI22XL addgen4_A_I2509 (.Y(N723), .A0(N724), .A1(N694), .B0(N722), .B1(N695));
XNOR2X1 addgen4_A_I2510 (.Y(N726), .A(N7682), .B(N7807));
OAI22XL addgen4_A_I2511 (.Y(N725), .A0(N726), .A1(N694), .B0(N724), .B1(N695));
XNOR2X1 addgen4_A_I2512 (.Y(N728), .A(N7683), .B(N7807));
OAI22XL addgen4_A_I2513 (.Y(N727), .A0(N728), .A1(N694), .B0(N726), .B1(N695));
XNOR2X1 addgen4_A_I2514 (.Y(N730), .A(N7684), .B(N7807));
OAI22XL addgen4_A_I2515 (.Y(N729), .A0(N730), .A1(N694), .B0(N728), .B1(N695));
XNOR2X1 addgen4_A_I2516 (.Y(N732), .A(N7685), .B(N7807));
OAI22XL addgen4_A_I2517 (.Y(N731), .A0(N732), .A1(N694), .B0(N730), .B1(N695));
XNOR2X1 addgen4_A_I2518 (.Y(N734), .A(N7686), .B(N7807));
OAI22XL addgen4_A_I2519 (.Y(N733), .A0(N734), .A1(N694), .B0(N732), .B1(N695));
XNOR2X1 addgen4_A_I2520 (.Y(N736), .A(N7687), .B(N7807));
OAI22XL addgen4_A_I2521 (.Y(N735), .A0(N736), .A1(N694), .B0(N734), .B1(N695));
XNOR2X1 addgen4_A_I2522 (.Y(N738), .A(N7688), .B(N7807));
OAI22XL addgen4_A_I2523 (.Y(N737), .A0(N738), .A1(N694), .B0(N736), .B1(N695));
XNOR2X1 addgen4_A_I2524 (.Y(N740), .A(N7689), .B(N7807));
OAI22XL addgen4_A_I2525 (.Y(N739), .A0(N740), .A1(N694), .B0(N738), .B1(N695));
XNOR2X1 addgen4_A_I2526 (.Y(N742), .A(N7690), .B(N7807));
OAI22XL addgen4_A_I2527 (.Y(N741), .A0(N742), .A1(N694), .B0(N740), .B1(N695));
XNOR2X1 addgen4_A_I2528 (.Y(N744), .A(N7691), .B(N7807));
OAI22XL addgen4_A_I2529 (.Y(N743), .A0(N744), .A1(N694), .B0(N742), .B1(N695));
XNOR2X1 addgen4_A_I2530 (.Y(N746), .A(N7692), .B(N7807));
OAI22XL addgen4_A_I2531 (.Y(N745), .A0(N746), .A1(N694), .B0(N744), .B1(N695));
INVXL addgen4_A_I2532 (.Y(N748), .A(N7807));
OAI22XL addgen4_A_I2533 (.Y(N747), .A0(N748), .A1(N694), .B0(N746), .B1(N695));
MXI2XL inst_cellmath__24_0_I273 (.Y(N749), .A(N695), .B(N694), .S0(N748));
XNOR2X1 enc3_A_I2534 (.Y(N758), .A(inst_cellmath__24_0_in0[12]), .B(inst_cellmath__24_0_in0[11]));
XOR2XL enc3_A_I2535 (.Y(N4872), .A(inst_cellmath__24_0_in0[13]), .B(inst_cellmath__24_0_in0[11]));
NAND2X2 enc3_A_I2537 (.Y(N759), .A(N4872), .B(N758));
INVX1 inst_cellmath__24_0_I3327 (.Y(N7829), .A(inst_cellmath__24_0_in0[13]));
NAND2XL inst_cellmath__24_0_I279 (.Y(N763), .A(inst_cellmath__24_0_in0[11]), .B(inst_cellmath__24_0_in0[12]));
AND2XL inst_cellmath__24_0_I280 (.Y(N764), .A(inst_cellmath__24_0_in0[13]), .B(N763));
XNOR2X1 addgen4_A_I2538 (.Y(N766), .A(N7670), .B(N7829));
OAI22XL addgen4_A_I2539 (.Y(N765), .A0(N766), .A1(N758), .B0(N7829), .B1(N759));
XNOR2X1 addgen4_A_I2540 (.Y(N768), .A(N7671), .B(N7829));
OAI22XL addgen4_A_I2541 (.Y(N767), .A0(N768), .A1(N758), .B0(N766), .B1(N759));
XNOR2X1 addgen4_A_I2542 (.Y(N770), .A(N7672), .B(N7829));
OAI22XL addgen4_A_I2543 (.Y(N769), .A0(N770), .A1(N758), .B0(N768), .B1(N759));
XNOR2X1 addgen4_A_I2544 (.Y(N772), .A(N7673), .B(N7829));
OAI22XL addgen4_A_I2545 (.Y(N771), .A0(N772), .A1(N758), .B0(N770), .B1(N759));
XNOR2X1 addgen4_A_I2546 (.Y(N774), .A(N7674), .B(N7829));
OAI22XL addgen4_A_I2547 (.Y(N773), .A0(N774), .A1(N758), .B0(N772), .B1(N759));
XNOR2X1 addgen4_A_I2548 (.Y(N776), .A(N7675), .B(N7829));
OAI22XL addgen4_A_I2549 (.Y(N775), .A0(N776), .A1(N758), .B0(N774), .B1(N759));
XNOR2X1 addgen4_A_I2550 (.Y(N778), .A(N7676), .B(N7829));
OAI22XL addgen4_A_I2551 (.Y(N777), .A0(N778), .A1(N758), .B0(N776), .B1(N759));
XNOR2X1 addgen4_A_I2552 (.Y(N780), .A(N7677), .B(N7829));
OAI22XL addgen4_A_I2553 (.Y(N779), .A0(N780), .A1(N758), .B0(N778), .B1(N759));
XNOR2X1 addgen4_A_I2554 (.Y(N782), .A(N7678), .B(N7829));
OAI22XL addgen4_A_I2555 (.Y(N781), .A0(N782), .A1(N758), .B0(N780), .B1(N759));
XNOR2X1 addgen4_A_I2556 (.Y(N784), .A(N7679), .B(N7829));
OAI22XL addgen4_A_I2557 (.Y(N783), .A0(N784), .A1(N758), .B0(N782), .B1(N759));
XNOR2X1 addgen4_A_I2558 (.Y(N786), .A(N7680), .B(N7829));
OAI22XL addgen4_A_I2559 (.Y(N785), .A0(N786), .A1(N758), .B0(N784), .B1(N759));
XNOR2X1 addgen4_A_I2560 (.Y(N788), .A(N7681), .B(N7829));
OAI22XL addgen4_A_I2561 (.Y(N787), .A0(N788), .A1(N758), .B0(N786), .B1(N759));
XNOR2X1 addgen4_A_I2562 (.Y(N790), .A(N7682), .B(N7829));
OAI22XL addgen4_A_I2563 (.Y(N789), .A0(N790), .A1(N758), .B0(N788), .B1(N759));
XNOR2X1 addgen4_A_I2564 (.Y(N792), .A(N7683), .B(N7829));
OAI22XL addgen4_A_I2565 (.Y(N791), .A0(N792), .A1(N758), .B0(N790), .B1(N759));
XNOR2X1 addgen4_A_I2566 (.Y(N794), .A(N7684), .B(N7829));
OAI22XL addgen4_A_I2567 (.Y(N793), .A0(N794), .A1(N758), .B0(N792), .B1(N759));
XNOR2X1 addgen4_A_I2568 (.Y(N796), .A(N7685), .B(N7829));
OAI22XL addgen4_A_I2569 (.Y(N795), .A0(N796), .A1(N758), .B0(N794), .B1(N759));
XNOR2X1 addgen4_A_I2570 (.Y(N798), .A(N7686), .B(N7829));
OAI22XL addgen4_A_I2571 (.Y(N797), .A0(N798), .A1(N758), .B0(N796), .B1(N759));
XNOR2X1 addgen4_A_I2572 (.Y(N800), .A(N7687), .B(N7829));
OAI22XL addgen4_A_I2573 (.Y(N799), .A0(N800), .A1(N758), .B0(N798), .B1(N759));
XNOR2X1 addgen4_A_I2574 (.Y(N802), .A(N7688), .B(N7829));
OAI22XL addgen4_A_I2575 (.Y(N801), .A0(N802), .A1(N758), .B0(N800), .B1(N759));
XNOR2X1 addgen4_A_I2576 (.Y(N804), .A(N7689), .B(N7829));
OAI22XL addgen4_A_I2577 (.Y(N803), .A0(N804), .A1(N758), .B0(N802), .B1(N759));
XNOR2X1 addgen4_A_I2578 (.Y(N806), .A(N7690), .B(N7829));
OAI22XL addgen4_A_I2579 (.Y(N805), .A0(N806), .A1(N758), .B0(N804), .B1(N759));
XNOR2X1 addgen4_A_I2580 (.Y(N808), .A(N7691), .B(N7829));
OAI22XL addgen4_A_I2581 (.Y(N807), .A0(N808), .A1(N758), .B0(N806), .B1(N759));
XNOR2X1 addgen4_A_I2582 (.Y(N810), .A(N7692), .B(N7829));
OAI22XL addgen4_A_I2583 (.Y(N809), .A0(N810), .A1(N758), .B0(N808), .B1(N759));
INVXL addgen4_A_I2584 (.Y(N812), .A(N7829));
OAI22XL addgen4_A_I2585 (.Y(N811), .A0(N812), .A1(N758), .B0(N810), .B1(N759));
MXI2XL inst_cellmath__24_0_I305 (.Y(N813), .A(N759), .B(N758), .S0(N812));
XNOR2X1 enc3_A_I2586 (.Y(N822), .A(inst_cellmath__24_0_in0[14]), .B(inst_cellmath__24_0_in0[13]));
XOR2XL enc3_A_I2587 (.Y(N5099), .A(inst_cellmath__24_0_in0[15]), .B(inst_cellmath__24_0_in0[13]));
NAND2X2 enc3_A_I2589 (.Y(N823), .A(N5099), .B(N822));
INVX1 inst_cellmath__24_0_I3339 (.Y(N7841), .A(inst_cellmath__24_0_in0[15]));
NAND2XL inst_cellmath__24_0_I311 (.Y(N827), .A(inst_cellmath__24_0_in0[13]), .B(inst_cellmath__24_0_in0[14]));
AND2XL inst_cellmath__24_0_I312 (.Y(N828), .A(inst_cellmath__24_0_in0[15]), .B(N827));
XNOR2X1 addgen4_A_I2590 (.Y(N830), .A(N7670), .B(N7841));
OAI22XL addgen4_A_I2591 (.Y(N829), .A0(N830), .A1(N822), .B0(N7841), .B1(N823));
XNOR2X1 addgen4_A_I2592 (.Y(N832), .A(N7671), .B(N7841));
OAI22XL addgen4_A_I2593 (.Y(N831), .A0(N832), .A1(N822), .B0(N830), .B1(N823));
XNOR2X1 addgen4_A_I2594 (.Y(N834), .A(N7672), .B(N7841));
OAI22XL addgen4_A_I2595 (.Y(N833), .A0(N834), .A1(N822), .B0(N832), .B1(N823));
XNOR2X1 addgen4_A_I2596 (.Y(N836), .A(N7673), .B(N7841));
OAI22XL addgen4_A_I2597 (.Y(N835), .A0(N836), .A1(N822), .B0(N834), .B1(N823));
XNOR2X1 addgen4_A_I2598 (.Y(N838), .A(N7674), .B(N7841));
OAI22XL addgen4_A_I2599 (.Y(N837), .A0(N838), .A1(N822), .B0(N836), .B1(N823));
XNOR2X1 addgen4_A_I2600 (.Y(N840), .A(N7675), .B(N7841));
OAI22XL addgen4_A_I2601 (.Y(N839), .A0(N840), .A1(N822), .B0(N838), .B1(N823));
XNOR2X1 addgen4_A_I2602 (.Y(N842), .A(N7676), .B(N7841));
OAI22XL addgen4_A_I2603 (.Y(N841), .A0(N842), .A1(N822), .B0(N840), .B1(N823));
XNOR2X1 addgen4_A_I2604 (.Y(N844), .A(N7677), .B(N7841));
OAI22XL addgen4_A_I2605 (.Y(N843), .A0(N844), .A1(N822), .B0(N842), .B1(N823));
XNOR2X1 addgen4_A_I2606 (.Y(N846), .A(N7678), .B(N7841));
OAI22XL addgen4_A_I2607 (.Y(N845), .A0(N846), .A1(N822), .B0(N844), .B1(N823));
XNOR2X1 addgen4_A_I2608 (.Y(N848), .A(N7679), .B(N7841));
OAI22XL addgen4_A_I2609 (.Y(N847), .A0(N848), .A1(N822), .B0(N846), .B1(N823));
XNOR2X1 addgen4_A_I2610 (.Y(N850), .A(N7680), .B(N7841));
OAI22XL addgen4_A_I2611 (.Y(N849), .A0(N850), .A1(N822), .B0(N848), .B1(N823));
XNOR2X1 addgen4_A_I2612 (.Y(N852), .A(N7681), .B(N7841));
OAI22XL addgen4_A_I2613 (.Y(N851), .A0(N852), .A1(N822), .B0(N850), .B1(N823));
XNOR2X1 addgen4_A_I2614 (.Y(N854), .A(N7682), .B(N7841));
OAI22XL addgen4_A_I2615 (.Y(N853), .A0(N854), .A1(N822), .B0(N852), .B1(N823));
XNOR2X1 addgen4_A_I2616 (.Y(N856), .A(N7683), .B(N7841));
OAI22XL addgen4_A_I2617 (.Y(N855), .A0(N856), .A1(N822), .B0(N854), .B1(N823));
XNOR2X1 addgen4_A_I2618 (.Y(N858), .A(N7684), .B(N7841));
OAI22XL addgen4_A_I2619 (.Y(N857), .A0(N858), .A1(N822), .B0(N856), .B1(N823));
XNOR2X1 addgen4_A_I2620 (.Y(N860), .A(N7685), .B(N7841));
OAI22XL addgen4_A_I2621 (.Y(N859), .A0(N860), .A1(N822), .B0(N858), .B1(N823));
XNOR2X1 addgen4_A_I2622 (.Y(N862), .A(N7686), .B(N7841));
OAI22XL addgen4_A_I2623 (.Y(N861), .A0(N862), .A1(N822), .B0(N860), .B1(N823));
XNOR2X1 addgen4_A_I2624 (.Y(N864), .A(N7687), .B(N7841));
OAI22XL addgen4_A_I2625 (.Y(N863), .A0(N864), .A1(N822), .B0(N862), .B1(N823));
XNOR2X1 addgen4_A_I2626 (.Y(N866), .A(N7688), .B(N7841));
OAI22XL addgen4_A_I2627 (.Y(N865), .A0(N866), .A1(N822), .B0(N864), .B1(N823));
XNOR2X1 addgen4_A_I2628 (.Y(N868), .A(N7689), .B(N7841));
OAI22XL addgen4_A_I2629 (.Y(N867), .A0(N868), .A1(N822), .B0(N866), .B1(N823));
XNOR2X1 addgen4_A_I2630 (.Y(N870), .A(N7690), .B(N7841));
OAI22XL addgen4_A_I2631 (.Y(N869), .A0(N870), .A1(N822), .B0(N868), .B1(N823));
XNOR2X1 addgen4_A_I2632 (.Y(N872), .A(N7691), .B(N7841));
OAI22XL addgen4_A_I2633 (.Y(N871), .A0(N872), .A1(N822), .B0(N870), .B1(N823));
XNOR2X1 addgen4_A_I2634 (.Y(N874), .A(N7692), .B(N7841));
OAI22XL addgen4_A_I2635 (.Y(N873), .A0(N874), .A1(N822), .B0(N872), .B1(N823));
INVXL addgen4_A_I2636 (.Y(N876), .A(N7841));
OAI22XL addgen4_A_I2637 (.Y(N875), .A0(N876), .A1(N822), .B0(N874), .B1(N823));
MXI2XL inst_cellmath__24_0_I337 (.Y(N877), .A(N823), .B(N822), .S0(N876));
XNOR2X1 enc3_A_I2638 (.Y(N886), .A(inst_cellmath__24_0_in0[16]), .B(inst_cellmath__24_0_in0[15]));
XOR2XL enc3_A_I2639 (.Y(N5326), .A(inst_cellmath__24_0_in0[17]), .B(inst_cellmath__24_0_in0[15]));
NAND2X2 enc3_A_I2641 (.Y(N887), .A(N5326), .B(N886));
INVX1 inst_cellmath__24_0_I3361 (.Y(N7863), .A(inst_cellmath__24_0_in0[17]));
NAND2XL inst_cellmath__24_0_I343 (.Y(N891), .A(inst_cellmath__24_0_in0[15]), .B(inst_cellmath__24_0_in0[16]));
AND2XL inst_cellmath__24_0_I344 (.Y(N892), .A(inst_cellmath__24_0_in0[17]), .B(N891));
XNOR2X1 addgen4_A_I2642 (.Y(N894), .A(N7670), .B(N7863));
OAI22XL addgen4_A_I2643 (.Y(N893), .A0(N894), .A1(N886), .B0(N7863), .B1(N887));
XNOR2X1 addgen4_A_I2644 (.Y(N896), .A(N7671), .B(N7863));
OAI22XL addgen4_A_I2645 (.Y(N895), .A0(N896), .A1(N886), .B0(N894), .B1(N887));
XNOR2X1 addgen4_A_I2646 (.Y(N898), .A(N7672), .B(N7863));
OAI22XL addgen4_A_I2647 (.Y(N897), .A0(N898), .A1(N886), .B0(N896), .B1(N887));
XNOR2X1 addgen4_A_I2648 (.Y(N900), .A(N7673), .B(N7863));
OAI22XL addgen4_A_I2649 (.Y(N899), .A0(N900), .A1(N886), .B0(N898), .B1(N887));
XNOR2X1 addgen4_A_I2650 (.Y(N902), .A(N7674), .B(N7863));
OAI22XL addgen4_A_I2651 (.Y(N901), .A0(N902), .A1(N886), .B0(N900), .B1(N887));
XNOR2X1 addgen4_A_I2652 (.Y(N904), .A(N7675), .B(N7863));
OAI22XL addgen4_A_I2653 (.Y(N903), .A0(N904), .A1(N886), .B0(N902), .B1(N887));
XNOR2X1 addgen4_A_I2654 (.Y(N906), .A(N7676), .B(N7863));
OAI22XL addgen4_A_I2655 (.Y(N905), .A0(N906), .A1(N886), .B0(N904), .B1(N887));
XNOR2X1 addgen4_A_I2656 (.Y(N908), .A(N7677), .B(N7863));
OAI22XL addgen4_A_I2657 (.Y(N907), .A0(N908), .A1(N886), .B0(N906), .B1(N887));
XNOR2X1 addgen4_A_I2658 (.Y(N910), .A(N7678), .B(N7863));
OAI22XL addgen4_A_I2659 (.Y(N909), .A0(N910), .A1(N886), .B0(N908), .B1(N887));
XNOR2X1 addgen4_A_I2660 (.Y(N912), .A(N7679), .B(N7863));
OAI22XL addgen4_A_I2661 (.Y(N911), .A0(N912), .A1(N886), .B0(N910), .B1(N887));
XNOR2X1 addgen4_A_I2662 (.Y(N914), .A(N7680), .B(N7863));
OAI22XL addgen4_A_I2663 (.Y(N913), .A0(N914), .A1(N886), .B0(N912), .B1(N887));
XNOR2X1 addgen4_A_I2664 (.Y(N916), .A(N7681), .B(N7863));
OAI22XL addgen4_A_I2665 (.Y(N915), .A0(N916), .A1(N886), .B0(N914), .B1(N887));
XNOR2X1 addgen4_A_I2666 (.Y(N918), .A(N7682), .B(N7863));
OAI22XL addgen4_A_I2667 (.Y(N917), .A0(N918), .A1(N886), .B0(N916), .B1(N887));
XNOR2X1 addgen4_A_I2668 (.Y(N920), .A(N7683), .B(N7863));
OAI22XL addgen4_A_I2669 (.Y(N919), .A0(N920), .A1(N886), .B0(N918), .B1(N887));
XNOR2X1 addgen4_A_I2670 (.Y(N922), .A(N7684), .B(N7863));
OAI22XL addgen4_A_I2671 (.Y(N921), .A0(N922), .A1(N886), .B0(N920), .B1(N887));
XNOR2X1 addgen4_A_I2672 (.Y(N924), .A(N7685), .B(N7863));
OAI22XL addgen4_A_I2673 (.Y(N923), .A0(N924), .A1(N886), .B0(N922), .B1(N887));
XNOR2X1 addgen4_A_I2674 (.Y(N926), .A(N7686), .B(N7863));
OAI22XL addgen4_A_I2675 (.Y(N925), .A0(N926), .A1(N886), .B0(N924), .B1(N887));
XNOR2X1 addgen4_A_I2676 (.Y(N928), .A(N7687), .B(N7863));
OAI22XL addgen4_A_I2677 (.Y(N927), .A0(N928), .A1(N886), .B0(N926), .B1(N887));
XNOR2X1 addgen4_A_I2678 (.Y(N930), .A(N7688), .B(N7863));
OAI22XL addgen4_A_I2679 (.Y(N929), .A0(N930), .A1(N886), .B0(N928), .B1(N887));
XNOR2X1 addgen4_A_I2680 (.Y(N932), .A(N7689), .B(N7863));
OAI22XL addgen4_A_I2681 (.Y(N931), .A0(N932), .A1(N886), .B0(N930), .B1(N887));
XNOR2X1 addgen4_A_I2682 (.Y(N934), .A(N7690), .B(N7863));
OAI22XL addgen4_A_I2683 (.Y(N933), .A0(N934), .A1(N886), .B0(N932), .B1(N887));
XNOR2X1 addgen4_A_I2684 (.Y(N936), .A(N7691), .B(N7863));
OAI22XL addgen4_A_I2685 (.Y(N935), .A0(N936), .A1(N886), .B0(N934), .B1(N887));
XNOR2X1 addgen4_A_I2686 (.Y(N938), .A(N7692), .B(N7863));
OAI22XL addgen4_A_I2687 (.Y(N937), .A0(N938), .A1(N886), .B0(N936), .B1(N887));
INVXL addgen4_A_I2688 (.Y(N940), .A(N7863));
OAI22XL addgen4_A_I2689 (.Y(N939), .A0(N940), .A1(N886), .B0(N938), .B1(N887));
MXI2XL inst_cellmath__24_0_I369 (.Y(N941), .A(N887), .B(N886), .S0(N940));
XNOR2X1 enc3_A_I2690 (.Y(N950), .A(inst_cellmath__24_0_in0[18]), .B(inst_cellmath__24_0_in0[17]));
XOR2XL enc3_A_I2691 (.Y(N5553), .A(inst_cellmath__24_0_in0[19]), .B(inst_cellmath__24_0_in0[17]));
NAND2X1 inst_cellmath__24_0_I3531 (.Y(N7874), .A(N5553), .B(N950));
INVXL inst_cellmath__24_0_I3373 (.Y(N7875), .A(inst_cellmath__24_0_in0[19]));
NAND2XL inst_cellmath__24_0_I375 (.Y(N955), .A(inst_cellmath__24_0_in0[17]), .B(inst_cellmath__24_0_in0[18]));
AND2XL inst_cellmath__24_0_I376 (.Y(N956), .A(inst_cellmath__24_0_in0[19]), .B(N955));
XNOR2X1 addgen4_A_I2694 (.Y(N958), .A(N7670), .B(N7875));
OAI22XL addgen4_A_I2695 (.Y(N957), .A0(N958), .A1(N950), .B0(N7875), .B1(N7874));
XNOR2X1 addgen4_A_I2696 (.Y(N960), .A(N7671), .B(N7875));
OAI22XL addgen4_A_I2697 (.Y(N959), .A0(N960), .A1(N950), .B0(N958), .B1(N7874));
XNOR2X1 addgen4_A_I2698 (.Y(N962), .A(N7672), .B(N7875));
OAI22XL addgen4_A_I2699 (.Y(N961), .A0(N962), .A1(N950), .B0(N960), .B1(N7874));
XNOR2X1 addgen4_A_I2700 (.Y(N964), .A(N7673), .B(N7875));
OAI22XL addgen4_A_I2701 (.Y(N963), .A0(N964), .A1(N950), .B0(N962), .B1(N7874));
XNOR2X1 addgen4_A_I2702 (.Y(N966), .A(N7674), .B(N7875));
OAI22XL addgen4_A_I2703 (.Y(N965), .A0(N966), .A1(N950), .B0(N964), .B1(N7874));
XNOR2X1 addgen4_A_I2704 (.Y(N968), .A(N7675), .B(N7875));
OAI22XL addgen4_A_I2705 (.Y(N967), .A0(N968), .A1(N950), .B0(N966), .B1(N7874));
XNOR2X1 addgen4_A_I2706 (.Y(N970), .A(N7676), .B(N7875));
OAI22XL addgen4_A_I2707 (.Y(N969), .A0(N970), .A1(N950), .B0(N968), .B1(N7874));
XNOR2X1 addgen4_A_I2708 (.Y(N972), .A(N7677), .B(N7875));
OAI22XL addgen4_A_I2709 (.Y(N971), .A0(N972), .A1(N950), .B0(N970), .B1(N7874));
XNOR2X1 addgen4_A_I2710 (.Y(N974), .A(N7678), .B(N7875));
OAI22XL addgen4_A_I2711 (.Y(N973), .A0(N974), .A1(N950), .B0(N972), .B1(N7874));
XNOR2X1 addgen4_A_I2712 (.Y(N976), .A(N7679), .B(N7875));
OAI22XL addgen4_A_I2713 (.Y(N975), .A0(N976), .A1(N950), .B0(N974), .B1(N7874));
XNOR2X1 addgen4_A_I2714 (.Y(N978), .A(N7680), .B(N7875));
OAI22XL addgen4_A_I2715 (.Y(N977), .A0(N978), .A1(N950), .B0(N976), .B1(N7874));
XNOR2X1 addgen4_A_I2716 (.Y(N980), .A(N7681), .B(N7875));
OAI22XL addgen4_A_I2717 (.Y(N979), .A0(N980), .A1(N950), .B0(N978), .B1(N7874));
XNOR2X1 addgen4_A_I2718 (.Y(N982), .A(N7682), .B(N7875));
OAI22XL addgen4_A_I2719 (.Y(N981), .A0(N982), .A1(N950), .B0(N980), .B1(N7874));
XNOR2X1 addgen4_A_I2720 (.Y(N984), .A(N7683), .B(N7875));
OAI22XL addgen4_A_I2721 (.Y(N983), .A0(N984), .A1(N950), .B0(N982), .B1(N7874));
XNOR2X1 addgen4_A_I2722 (.Y(N986), .A(N7684), .B(N7875));
OAI22XL addgen4_A_I2723 (.Y(N985), .A0(N986), .A1(N950), .B0(N984), .B1(N7874));
XNOR2X1 addgen4_A_I2724 (.Y(N988), .A(N7685), .B(N7875));
OAI22XL addgen4_A_I2725 (.Y(N987), .A0(N988), .A1(N950), .B0(N986), .B1(N7874));
XNOR2X1 addgen4_A_I2726 (.Y(N990), .A(N7686), .B(N7875));
OAI22XL addgen4_A_I2727 (.Y(N989), .A0(N990), .A1(N950), .B0(N988), .B1(N7874));
XNOR2X1 addgen4_A_I2728 (.Y(N992), .A(N7687), .B(N7875));
OAI22XL addgen4_A_I2729 (.Y(N991), .A0(N992), .A1(N950), .B0(N990), .B1(N7874));
XNOR2X1 addgen4_A_I2730 (.Y(N994), .A(N7688), .B(N7875));
OAI22XL addgen4_A_I2731 (.Y(N993), .A0(N994), .A1(N950), .B0(N992), .B1(N7874));
XNOR2X1 addgen4_A_I2732 (.Y(N996), .A(N7689), .B(N7875));
OAI22XL addgen4_A_I2733 (.Y(N995), .A0(N996), .A1(N950), .B0(N994), .B1(N7874));
XNOR2X1 addgen4_A_I2734 (.Y(N998), .A(N7690), .B(N7875));
OAI22XL addgen4_A_I2735 (.Y(N997), .A0(N998), .A1(N950), .B0(N996), .B1(N7874));
XNOR2X1 addgen4_A_I2736 (.Y(N1000), .A(N7691), .B(N7875));
OAI22XL addgen4_A_I2737 (.Y(N999), .A0(N1000), .A1(N950), .B0(N998), .B1(N7874));
XNOR2X1 addgen4_A_I2738 (.Y(N1002), .A(N7692), .B(N7875));
OAI22XL addgen4_A_I2739 (.Y(N1001), .A0(N1002), .A1(N950), .B0(N1000), .B1(N7874));
INVXL addgen4_A_I2740 (.Y(N1004), .A(N7875));
OAI22XL addgen4_A_I2741 (.Y(N1003), .A0(N1004), .A1(N950), .B0(N1002), .B1(N7874));
MXI2XL inst_cellmath__24_0_I401 (.Y(N1005), .A(N7874), .B(N950), .S0(N1004));
XNOR2X1 enc3_A_I2742 (.Y(N1014), .A(inst_cellmath__24_0_in0[20]), .B(inst_cellmath__24_0_in0[19]));
XOR2XL enc3_A_I2743 (.Y(N5780), .A(inst_cellmath__24_0_in0[21]), .B(inst_cellmath__24_0_in0[19]));
NAND2X1 inst_cellmath__24_0_I3533 (.Y(N7886), .A(N5780), .B(N1014));
INVXL inst_cellmath__24_0_I3385 (.Y(N7887), .A(inst_cellmath__24_0_in0[21]));
NAND2XL inst_cellmath__24_0_I407 (.Y(N1019), .A(inst_cellmath__24_0_in0[19]), .B(inst_cellmath__24_0_in0[20]));
AND2XL inst_cellmath__24_0_I408 (.Y(N1020), .A(inst_cellmath__24_0_in0[21]), .B(N1019));
XNOR2X1 addgen4_A_I2746 (.Y(N1022), .A(N7670), .B(N7887));
OAI22XL addgen4_A_I2747 (.Y(N1021), .A0(N1022), .A1(N1014), .B0(N7887), .B1(N7886));
XNOR2X1 addgen4_A_I2748 (.Y(N1024), .A(N7671), .B(N7887));
OAI22XL addgen4_A_I2749 (.Y(N1023), .A0(N1024), .A1(N1014), .B0(N1022), .B1(N7886));
XNOR2X1 addgen4_A_I2750 (.Y(N1026), .A(N7672), .B(N7887));
OAI22XL addgen4_A_I2751 (.Y(N1025), .A0(N1026), .A1(N1014), .B0(N1024), .B1(N7886));
XNOR2X1 addgen4_A_I2752 (.Y(N1028), .A(N7673), .B(N7887));
OAI22XL addgen4_A_I2753 (.Y(N1027), .A0(N1028), .A1(N1014), .B0(N1026), .B1(N7886));
XNOR2X1 addgen4_A_I2754 (.Y(N1030), .A(N7674), .B(N7887));
OAI22XL addgen4_A_I2755 (.Y(N1029), .A0(N1030), .A1(N1014), .B0(N1028), .B1(N7886));
XNOR2X1 addgen4_A_I2756 (.Y(N1032), .A(N7675), .B(N7887));
OAI22XL addgen4_A_I2757 (.Y(N1031), .A0(N1032), .A1(N1014), .B0(N1030), .B1(N7886));
XNOR2X1 addgen4_A_I2758 (.Y(N1034), .A(N7676), .B(N7887));
OAI22XL addgen4_A_I2759 (.Y(N1033), .A0(N1034), .A1(N1014), .B0(N1032), .B1(N7886));
XNOR2X1 addgen4_A_I2760 (.Y(N1036), .A(N7677), .B(N7887));
OAI22XL addgen4_A_I2761 (.Y(N1035), .A0(N1036), .A1(N1014), .B0(N1034), .B1(N7886));
XNOR2X1 addgen4_A_I2762 (.Y(N1038), .A(N7678), .B(N7887));
OAI22XL addgen4_A_I2763 (.Y(N1037), .A0(N1038), .A1(N1014), .B0(N1036), .B1(N7886));
XNOR2X1 addgen4_A_I2764 (.Y(N1040), .A(N7679), .B(N7887));
OAI22XL addgen4_A_I2765 (.Y(N1039), .A0(N1040), .A1(N1014), .B0(N1038), .B1(N7886));
XNOR2X1 addgen4_A_I2766 (.Y(N1042), .A(N7680), .B(N7887));
OAI22XL addgen4_A_I2767 (.Y(N1041), .A0(N1042), .A1(N1014), .B0(N1040), .B1(N7886));
XNOR2X1 addgen4_A_I2768 (.Y(N1044), .A(N7681), .B(N7887));
OAI22XL addgen4_A_I2769 (.Y(N1043), .A0(N1044), .A1(N1014), .B0(N1042), .B1(N7886));
XNOR2X1 addgen4_A_I2770 (.Y(N1046), .A(N7682), .B(N7887));
OAI22XL addgen4_A_I2771 (.Y(N1045), .A0(N1046), .A1(N1014), .B0(N1044), .B1(N7886));
XNOR2X1 addgen4_A_I2772 (.Y(N1048), .A(N7683), .B(N7887));
OAI22XL addgen4_A_I2773 (.Y(N1047), .A0(N1048), .A1(N1014), .B0(N1046), .B1(N7886));
XNOR2X1 addgen4_A_I2774 (.Y(N1050), .A(N7684), .B(N7887));
OAI22XL addgen4_A_I2775 (.Y(N1049), .A0(N1050), .A1(N1014), .B0(N1048), .B1(N7886));
XNOR2X1 addgen4_A_I2776 (.Y(N1052), .A(N7685), .B(N7887));
OAI22XL addgen4_A_I2777 (.Y(N1051), .A0(N1052), .A1(N1014), .B0(N1050), .B1(N7886));
XNOR2X1 addgen4_A_I2778 (.Y(N1054), .A(N7686), .B(N7887));
OAI22XL addgen4_A_I2779 (.Y(N1053), .A0(N1054), .A1(N1014), .B0(N1052), .B1(N7886));
XNOR2X1 addgen4_A_I2780 (.Y(N1056), .A(N7687), .B(N7887));
OAI22XL addgen4_A_I2781 (.Y(N1055), .A0(N1056), .A1(N1014), .B0(N1054), .B1(N7886));
XNOR2X1 addgen4_A_I2782 (.Y(N1058), .A(N7688), .B(N7887));
OAI22XL addgen4_A_I2783 (.Y(N1057), .A0(N1058), .A1(N1014), .B0(N1056), .B1(N7886));
XNOR2X1 addgen4_A_I2784 (.Y(N1060), .A(N7689), .B(N7887));
OAI22XL addgen4_A_I2785 (.Y(N1059), .A0(N1060), .A1(N1014), .B0(N1058), .B1(N7886));
XNOR2X1 addgen4_A_I2786 (.Y(N1062), .A(N7690), .B(N7887));
OAI22XL addgen4_A_I2787 (.Y(N1061), .A0(N1062), .A1(N1014), .B0(N1060), .B1(N7886));
XNOR2X1 addgen4_A_I2788 (.Y(N1064), .A(N7691), .B(N7887));
OAI22XL addgen4_A_I2789 (.Y(N1063), .A0(N1064), .A1(N1014), .B0(N1062), .B1(N7886));
XNOR2X1 addgen4_A_I2790 (.Y(N1066), .A(N7692), .B(N7887));
OAI22XL addgen4_A_I2791 (.Y(N1065), .A0(N1066), .A1(N1014), .B0(N1064), .B1(N7886));
INVXL addgen4_A_I2792 (.Y(N1068), .A(N7887));
OAI22XL addgen4_A_I2793 (.Y(N1067), .A0(N1068), .A1(N1014), .B0(N1066), .B1(N7886));
MXI2XL inst_cellmath__24_0_I433 (.Y(N1069), .A(N7886), .B(N1014), .S0(N1068));
XNOR2X1 inst_cellmath__24_0_I2794 (.Y(N1078), .A(inst_cellmath__24_0_in0[22]), .B(inst_cellmath__24_0_in0[21]));
OR2XL inst_cellmath__24_0_I3534 (.Y(N7907), .A(inst_cellmath__24_0_in0[22]), .B(inst_cellmath__24_0_in0[21]));
NAND2XL inst_cellmath__24_0_I439 (.Y(N1084), .A(inst_cellmath__24_0_in0[21]), .B(inst_cellmath__24_0_in0[22]));
INVXL addgen4_A_I2796 (.Y(N1093), .A(N7670));
OAI21XL addgen4_A_I2797 (.Y(N1092), .A0(N1078), .A1(N1093), .B0(N7907));
INVXL addgen4_A_I2798 (.Y(N1095), .A(N7671));
OAI22XL addgen4_A_I2799 (.Y(N1094), .A0(N1095), .A1(N1078), .B0(N1093), .B1(N7907));
INVXL addgen4_A_I2800 (.Y(N1097), .A(N7672));
OAI22XL addgen4_A_I2801 (.Y(N1096), .A0(N1097), .A1(N1078), .B0(N1095), .B1(N7907));
INVXL addgen4_A_I2802 (.Y(N1099), .A(N7673));
OAI22XL addgen4_A_I2803 (.Y(N1098), .A0(N1099), .A1(N1078), .B0(N1097), .B1(N7907));
INVXL addgen4_A_I2804 (.Y(N1101), .A(N7674));
OAI22XL addgen4_A_I2805 (.Y(N1100), .A0(N1101), .A1(N1078), .B0(N1099), .B1(N7907));
INVXL addgen4_A_I2806 (.Y(N1103), .A(N7675));
OAI22XL addgen4_A_I2807 (.Y(N1102), .A0(N1103), .A1(N1078), .B0(N1101), .B1(N7907));
INVXL addgen4_A_I2808 (.Y(N1105), .A(N7676));
OAI22XL addgen4_A_I2809 (.Y(N1104), .A0(N1105), .A1(N1078), .B0(N1103), .B1(N7907));
INVXL addgen4_A_I2810 (.Y(N1107), .A(N7677));
OAI22XL addgen4_A_I2811 (.Y(N1106), .A0(N1107), .A1(N1078), .B0(N1105), .B1(N7907));
INVXL addgen4_A_I2812 (.Y(N1109), .A(N7678));
OAI22XL addgen4_A_I2813 (.Y(N1108), .A0(N1109), .A1(N1078), .B0(N1107), .B1(N7907));
INVXL addgen4_A_I2814 (.Y(N1111), .A(N7679));
OAI22XL addgen4_A_I2815 (.Y(N1110), .A0(N1111), .A1(N1078), .B0(N1109), .B1(N7907));
INVXL addgen4_A_I2816 (.Y(N1113), .A(N7680));
OAI22XL addgen4_A_I2817 (.Y(N1112), .A0(N1113), .A1(N1078), .B0(N1111), .B1(N7907));
INVXL addgen4_A_I2818 (.Y(N1115), .A(N7681));
OAI22XL addgen4_A_I2819 (.Y(N1114), .A0(N1115), .A1(N1078), .B0(N1113), .B1(N7907));
INVXL addgen4_A_I2820 (.Y(N1117), .A(N7682));
OAI22XL addgen4_A_I2821 (.Y(N1116), .A0(N1117), .A1(N1078), .B0(N1115), .B1(N7907));
INVXL addgen4_A_I2822 (.Y(N1119), .A(N7683));
OAI22XL addgen4_A_I2823 (.Y(N1118), .A0(N1119), .A1(N1078), .B0(N1117), .B1(N7907));
INVXL addgen4_A_I2824 (.Y(N1121), .A(N7684));
OAI22XL addgen4_A_I2825 (.Y(N1120), .A0(N1121), .A1(N1078), .B0(N1119), .B1(N7907));
INVXL addgen4_A_I2826 (.Y(N1123), .A(N7685));
OAI22XL addgen4_A_I2827 (.Y(N1122), .A0(N1123), .A1(N1078), .B0(N1121), .B1(N7907));
INVXL addgen4_A_I2828 (.Y(N1125), .A(N7686));
OAI22XL addgen4_A_I2829 (.Y(N1124), .A0(N1125), .A1(N1078), .B0(N1123), .B1(N7907));
INVXL addgen4_A_I2830 (.Y(N1127), .A(N7687));
OAI22XL addgen4_A_I2831 (.Y(N1126), .A0(N1127), .A1(N1078), .B0(N1125), .B1(N7907));
INVXL addgen4_A_I2832 (.Y(N1129), .A(N7688));
OAI22XL addgen4_A_I2833 (.Y(N1128), .A0(N1129), .A1(N1078), .B0(N1127), .B1(N7907));
INVXL addgen4_A_I2834 (.Y(N1131), .A(N7689));
OAI22XL addgen4_A_I2835 (.Y(N1130), .A0(N1131), .A1(N1078), .B0(N1129), .B1(N7907));
INVXL addgen4_A_I2836 (.Y(N1133), .A(N7690));
OAI22XL addgen4_A_I2837 (.Y(N1132), .A0(N1133), .A1(N1078), .B0(N1131), .B1(N7907));
INVXL addgen4_A_I2838 (.Y(N1135), .A(N7691));
OAI22XL addgen4_A_I2839 (.Y(N1134), .A0(N1135), .A1(N1078), .B0(N1133), .B1(N7907));
INVXL addgen4_A_I2840 (.Y(N1137), .A(N7692));
OAI22XL addgen4_A_I2841 (.Y(N1136), .A0(N1137), .A1(N1078), .B0(N1135), .B1(N7907));
NOR2XL inst_cellmath__24_0_I464 (.Y(N1138), .A(N1137), .B(N7907));
INVXL inst_cellmath__24_0_I465 (.Y(N1140), .A(N1078));
NAND2XL inst_cellmath__24_0_I466 (.Y(N1144), .A(N1078), .B(N7907));
AO21XL inst_cellmath__24_0_I3147 (.Y(N1212), .A0(N372), .A1(N7696), .B0(N7697));
AO21XL inst_cellmath__24_0_I3148 (.Y(N1213), .A0(N438), .A1(N7718), .B0(N7719));
AO21XL inst_cellmath__24_0_I3149 (.Y(N1214), .A0(N502), .A1(N7740), .B0(N7741));
AO21XL inst_cellmath__24_0_I3150 (.Y(N1215), .A0(N566), .A1(N567), .B0(N7763));
AO21XL inst_cellmath__24_0_I3151 (.Y(N1216), .A0(N630), .A1(N631), .B0(N7785));
AO21XL inst_cellmath__24_0_I3152 (.Y(N1217), .A0(N694), .A1(N695), .B0(N7807));
AO21XL inst_cellmath__24_0_I3153 (.Y(N1218), .A0(N758), .A1(N759), .B0(N7829));
AO21XL inst_cellmath__24_0_I3154 (.Y(N1219), .A0(N822), .A1(N823), .B0(N7841));
AO21XL inst_cellmath__24_0_I3155 (.Y(N1220), .A0(N886), .A1(N887), .B0(N7863));
AO21XL inst_cellmath__24_0_I3156 (.Y(N1221), .A0(N950), .A1(N7874), .B0(N7875));
AO21XL inst_cellmath__24_0_I3157 (.Y(N1222), .A0(N1014), .A1(N7886), .B0(N7887));
ADDHX1 inst_cellmath__24_0_I510 (.CO(N1224), .S(N1223), .A(N444), .B(N385));
ADDHX1 inst_cellmath__24_0_I511 (.CO(N1226), .S(N1225), .A(N387), .B(N447));
ADDHX1 inst_cellmath__24_0_I512 (.CO(N1228), .S(N1227), .A(N508), .B(N389));
ADDFX1 inst_cellmath__24_0_I513 (.CO(N1230), .S(N1229), .A(N509), .B(N449), .CI(N1226));
ADDHX1 inst_cellmath__24_0_I514 (.CO(N1232), .S(N1231), .A(N391), .B(N451));
ADDFX1 inst_cellmath__24_0_I515 (.CO(N1234), .S(N1233), .A(N1228), .B(N511), .CI(N1231));
ADDHX1 inst_cellmath__24_0_I516 (.CO(N1236), .S(N1235), .A(N572), .B(N393));
ADDFX1 arith_dfa_A_I2842 (.CO(N1239), .S(N6216), .A(N513), .B(N453), .CI(N573));
ADDFX1 arith_dfa_A_I2843 (.CO(N1238), .S(N1237), .A(N1232), .B(N1235), .CI(N6216));
ADDHX1 inst_cellmath__24_0_I518 (.CO(N1241), .S(N1240), .A(N395), .B(N455));
ADDFX1 inst_cellmath__24_0_I519 (.CO(N1246), .S(N1245), .A(N575), .B(N515), .CI(N1236));
ADDFX1 inst_cellmath__24_0_I520 (.CO(N1248), .S(N1247), .A(N1239), .B(N1240), .CI(N1245));
ADDHX1 inst_cellmath__24_0_I521 (.CO(N1250), .S(N1249), .A(N636), .B(N397));
ADDFX1 inst_cellmath__24_0_I522 (.CO(N1252), .S(N1251), .A(N517), .B(N457), .CI(N577));
ADDFX1 arith_dfa_A_I2844 (.CO(N1255), .S(N6229), .A(N1241), .B(N637), .CI(N1249));
ADDFX1 arith_dfa_A_I2845 (.CO(N1254), .S(N1253), .A(N1246), .B(N1251), .CI(N6229));
ADDHX1 inst_cellmath__24_0_I524 (.CO(N1257), .S(N1256), .A(N399), .B(N459));
ADDFX1 inst_cellmath__24_0_I525 (.CO(N1259), .S(N1258), .A(N579), .B(N519), .CI(N639));
ADDFX1 inst_cellmath__24_0_I526 (.CO(N1264), .S(N1263), .A(N1256), .B(N1250), .CI(N1252));
ADDFX1 inst_cellmath__24_0_I527 (.CO(N1266), .S(N1265), .A(N1258), .B(N1255), .CI(N1263));
ADDHX1 inst_cellmath__24_0_I528 (.CO(N1268), .S(N1267), .A(N700), .B(N401));
ADDFX1 arith_dfa_A_I2846 (.CO(N1271), .S(N6242), .A(N521), .B(N461), .CI(N581));
ADDFX1 arith_dfa_A_I2847 (.CO(N1270), .S(N1269), .A(N1259), .B(N1267), .CI(N6242));
ADDFX1 inst_cellmath__24_0_I530 (.CO(N1276), .S(N1275), .A(N701), .B(N641), .CI(N1257));
ADDFX1 inst_cellmath__24_0_I531 (.CO(N1278), .S(N1277), .A(N1264), .B(N1275), .CI(N1269));
ADDHX1 inst_cellmath__24_0_I532 (.CO(N1280), .S(N1279), .A(N403), .B(N463));
ADDFX1 arith_dfa_A_I2848 (.CO(N1283), .S(N6255), .A(N583), .B(N523), .CI(N643));
ADDFX1 arith_dfa_A_I2849 (.CO(N1282), .S(N1281), .A(N1279), .B(N1271), .CI(N6255));
ADDFX1 inst_cellmath__24_0_I534 (.CO(N1288), .S(N1287), .A(N1268), .B(N703), .CI(N1276));
ADDFX1 inst_cellmath__24_0_I535 (.CO(N1290), .S(N1289), .A(N1287), .B(N1270), .CI(N1281));
ADDHX1 inst_cellmath__24_0_I536 (.CO(N1292), .S(N1291), .A(N764), .B(N405));
ADDFX1 inst_cellmath__24_0_I537 (.CO(N1294), .S(N1293), .A(N525), .B(N465), .CI(N585));
ADDFX1 arith_dfa_A_I2850 (.CO(N1297), .S(N6268), .A(N705), .B(N645), .CI(N765));
ADDFX1 arith_dfa_A_I2851 (.CO(N1296), .S(N1295), .A(N1291), .B(N1283), .CI(N6268));
ADDFX1 inst_cellmath__24_0_I539 (.CO(N1302), .S(N1301), .A(N1293), .B(N1280), .CI(N1288));
ADDFX1 inst_cellmath__24_0_I540 (.CO(N1304), .S(N1303), .A(N1295), .B(N1282), .CI(N1301));
ADDHX1 inst_cellmath__24_0_I541 (.CO(N1306), .S(N1305), .A(N407), .B(N467));
ADDFX1 inst_cellmath__24_0_I542 (.CO(N1308), .S(N1307), .A(N587), .B(N527), .CI(N647));
ADDFX1 inst_cellmath__24_0_I543 (.CO(N1313), .S(N1312), .A(N767), .B(N707), .CI(N1292));
ADDFX1 inst_cellmath__24_0_I544 (.CO(N1315), .S(N1314), .A(N1297), .B(N1305), .CI(N1294));
ADDFX1 inst_cellmath__24_0_I545 (.CO(N1320), .S(N1319), .A(N1312), .B(N1307), .CI(N1296));
ADDFX1 inst_cellmath__24_0_I546 (.CO(N1322), .S(N1321), .A(N1302), .B(N1314), .CI(N1319));
ADDHX1 inst_cellmath__24_0_I547 (.CO(N1324), .S(N1323), .A(N828), .B(N409));
ADDFX1 arith_dfa_A_I2852 (.CO(N1327), .S(N6281), .A(N529), .B(N469), .CI(N589));
ADDFX1 arith_dfa_A_I2853 (.CO(N1326), .S(N1325), .A(N1308), .B(N1323), .CI(N6281));
ADDFX1 arith_dfa_A_I2854 (.CO(N1330), .S(N6294), .A(N709), .B(N649), .CI(N769));
ADDFX1 arith_dfa_A_I2855 (.CO(N1329), .S(N1328), .A(N829), .B(N1306), .CI(N6294));
ADDFX1 inst_cellmath__24_0_I550 (.CO(N1335), .S(N1334), .A(N1315), .B(N1313), .CI(N1325));
ADDFX1 inst_cellmath__24_0_I551 (.CO(N1337), .S(N1336), .A(N1320), .B(N1328), .CI(N1334));
ADDHX1 inst_cellmath__24_0_I552 (.CO(N1339), .S(N1338), .A(N411), .B(N471));
ADDFX1 arith_dfa_A_I2856 (.CO(N1342), .S(N6307), .A(N591), .B(N531), .CI(N651));
ADDFX1 arith_dfa_A_I2857 (.CO(N1341), .S(N1340), .A(N1330), .B(N1327), .CI(N6307));
ADDFX1 arith_dfa_A_I2858 (.CO(N1345), .S(N6320), .A(N771), .B(N711), .CI(N831));
ADDFX1 arith_dfa_A_I2859 (.CO(N1344), .S(N1343), .A(N1324), .B(N1338), .CI(N6320));
ADDFX1 inst_cellmath__24_0_I555 (.CO(N1350), .S(N1349), .A(N1329), .B(N1326), .CI(N1340));
ADDFX1 inst_cellmath__24_0_I556 (.CO(N1352), .S(N1351), .A(N1335), .B(N1343), .CI(N1349));
ADDHX1 inst_cellmath__24_0_I557 (.CO(N1354), .S(N1353), .A(N892), .B(N413));
ADDFX1 inst_cellmath__24_0_I558 (.CO(N1356), .S(N1355), .A(N533), .B(N473), .CI(N593));
ADDFX1 arith_dfa_A_I2860 (.CO(N1359), .S(N6333), .A(N713), .B(N653), .CI(N773));
ADDFX1 arith_dfa_A_I2861 (.CO(N1358), .S(N1357), .A(N1345), .B(N1342), .CI(N6333));
ADDFX1 inst_cellmath__24_0_I560 (.CO(N1364), .S(N1363), .A(N833), .B(N893), .CI(N1339));
ADDFX1 inst_cellmath__24_0_I561 (.CO(N1366), .S(N1365), .A(N1355), .B(N1353), .CI(N1363));
ADDFX1 inst_cellmath__24_0_I562 (.CO(N1371), .S(N1370), .A(N1344), .B(N1341), .CI(N1365));
ADDFX1 inst_cellmath__24_0_I563 (.CO(N1373), .S(N1372), .A(N1350), .B(N1357), .CI(N1370));
ADDHX1 inst_cellmath__24_0_I564 (.CO(N1375), .S(N1374), .A(N415), .B(N475));
ADDFX1 inst_cellmath__24_0_I565 (.CO(N1377), .S(N1376), .A(N595), .B(N535), .CI(N655));
ADDFX1 arith_dfa_A_I2862 (.CO(N1380), .S(N6346), .A(N775), .B(N715), .CI(N835));
ADDFX1 arith_dfa_A_I2863 (.CO(N1379), .S(N1378), .A(N1356), .B(N1359), .CI(N6346));
ADDFX1 inst_cellmath__24_0_I567 (.CO(N1385), .S(N1384), .A(N1354), .B(N895), .CI(N1374));
ADDFX1 inst_cellmath__24_0_I568 (.CO(N1387), .S(N1386), .A(N1376), .B(N1364), .CI(N1384));
ADDFX1 inst_cellmath__24_0_I569 (.CO(N1392), .S(N1391), .A(N1366), .B(N1358), .CI(N1378));
ADDFX1 inst_cellmath__24_0_I570 (.CO(N1394), .S(N1393), .A(N1371), .B(N1386), .CI(N1391));
ADDHX1 inst_cellmath__24_0_I571 (.CO(N1396), .S(N1395), .A(N956), .B(N417));
ADDFX1 arith_dfa_A_I2864 (.CO(N1399), .S(N6359), .A(N477), .B(N597), .CI(N537));
ADDFX1 arith_dfa_A_I2865 (.CO(N1398), .S(N1397), .A(N1377), .B(N1380), .CI(N6359));
ADDFX1 arith_dfa_A_I2866 (.CO(N1402), .S(N6372), .A(N717), .B(N657), .CI(N777));
ADDFX1 arith_dfa_A_I2867 (.CO(N1401), .S(N1400), .A(N1375), .B(N1395), .CI(N6372));
ADDFX1 inst_cellmath__24_0_I574 (.CO(N1407), .S(N1406), .A(N897), .B(N837), .CI(N957));
ADDFX1 inst_cellmath__24_0_I575 (.CO(N1409), .S(N1408), .A(N1385), .B(N1406), .CI(N1379));
ADDFX1 arith_dfa_A_I2868 (.CO(N1412), .S(N6385), .A(N1397), .B(N1387), .CI(N1400));
ADDFX1 arith_dfa_A_I2869 (.CO(N1411), .S(N1410), .A(N1392), .B(N1408), .CI(N6385));
ADDHX1 inst_cellmath__24_0_I577 (.CO(N1414), .S(N1413), .A(N419), .B(N479));
ADDFX1 arith_dfa_A_I2870 (.CO(N1417), .S(N6398), .A(N599), .B(N539), .CI(N659));
ADDFX1 arith_dfa_A_I2871 (.CO(N1416), .S(N1415), .A(N1407), .B(N1399), .CI(N6398));
ADDFX1 arith_dfa_A_I2872 (.CO(N1420), .S(N6411), .A(N779), .B(N719), .CI(N839));
ADDFX1 arith_dfa_A_I2873 (.CO(N1419), .S(N1418), .A(N1413), .B(N1402), .CI(N6411));
ADDFX1 inst_cellmath__24_0_I580 (.CO(N1425), .S(N1424), .A(N959), .B(N899), .CI(N1396));
ADDFX1 inst_cellmath__24_0_I581 (.CO(N1427), .S(N1426), .A(N1398), .B(N1424), .CI(N1401));
ADDFX1 arith_dfa_A_I2874 (.CO(N1430), .S(N6424), .A(N1418), .B(N1415), .CI(N1409));
ADDFX1 arith_dfa_A_I2875 (.CO(N1429), .S(N1428), .A(N1426), .B(N1412), .CI(N6424));
ADDHX1 inst_cellmath__24_0_I583 (.CO(N1432), .S(N1431), .A(N1020), .B(N421));
ADDFX1 inst_cellmath__24_0_I584 (.CO(N1434), .S(N1433), .A(N541), .B(N481), .CI(N601));
ADDFX1 arith_dfa_A_I2876 (.CO(N1437), .S(N6437), .A(N721), .B(N661), .CI(N781));
ADDFX1 arith_dfa_A_I2877 (.CO(N1436), .S(N1435), .A(N1420), .B(N1417), .CI(N6437));
ADDFX1 arith_dfa_A_I2878 (.CO(N1440), .S(N6450), .A(N901), .B(N841), .CI(N961));
ADDFX1 arith_dfa_A_I2879 (.CO(N1439), .S(N1438), .A(N1414), .B(N1431), .CI(N6450));
ADDFX1 inst_cellmath__24_0_I587 (.CO(N1445), .S(N1444), .A(N1425), .B(N1021), .CI(N1433));
ADDFX1 inst_cellmath__24_0_I588 (.CO(N1447), .S(N1446), .A(N1419), .B(N1416), .CI(N1444));
ADDFX1 arith_dfa_A_I2880 (.CO(N1450), .S(N6463), .A(N1438), .B(N1435), .CI(N1427));
ADDFX1 arith_dfa_A_I2881 (.CO(N1449), .S(N1448), .A(N1446), .B(N1430), .CI(N6463));
ADDHX1 inst_cellmath__24_0_I590 (.CO(N1452), .S(N1451), .A(N423), .B(N483));
ADDFX1 inst_cellmath__24_0_I591 (.CO(N1454), .S(N1453), .A(N603), .B(N543), .CI(N663));
ADDFX1 arith_dfa_A_I2882 (.CO(N1457), .S(N6476), .A(N783), .B(N723), .CI(N843));
ADDFX1 arith_dfa_A_I2883 (.CO(N1456), .S(N1455), .A(N1434), .B(N1437), .CI(N6476));
ADDFX1 arith_dfa_A_I2884 (.CO(N1460), .S(N6489), .A(N963), .B(N903), .CI(N1023));
ADDFX1 arith_dfa_A_I2885 (.CO(N1459), .S(N1458), .A(N1451), .B(N1440), .CI(N6489));
ADDFX1 inst_cellmath__24_0_I594 (.CO(N1465), .S(N1464), .A(N1453), .B(N1432), .CI(N1445));
ADDFX1 inst_cellmath__24_0_I595 (.CO(N1467), .S(N1466), .A(N1439), .B(N1436), .CI(N1458));
ADDFX1 inst_cellmath__24_0_I596 (.CO(N1472), .S(N1471), .A(N1447), .B(N1455), .CI(N1464));
ADDFX1 inst_cellmath__24_0_I597 (.CO(N1474), .S(N1473), .A(N1450), .B(N1466), .CI(N1471));
ADDHX1 inst_cellmath__24_0_I598 (.CO(N1476), .S(N1475), .A(N1084), .B(N1092));
ADDFX1 arith_dfa_A_I2886 (.CO(N1479), .S(N6502), .A(N485), .B(N425), .CI(N545));
ADDFX1 arith_dfa_A_I2887 (.CO(N1478), .S(N1477), .A(N1454), .B(N1457), .CI(N6502));
ADDFX1 arith_dfa_A_I2888 (.CO(N1482), .S(N6515), .A(N665), .B(N605), .CI(N725));
ADDFX1 arith_dfa_A_I2889 (.CO(N1481), .S(N1480), .A(N1452), .B(N1460), .CI(N6515));
ADDFX1 inst_cellmath__24_0_I601 (.CO(N1487), .S(N1486), .A(N785), .B(N1025), .CI(N845));
ADDFX1 inst_cellmath__24_0_I602 (.CO(N1489), .S(N1488), .A(N965), .B(N905), .CI(N1475));
ADDFX1 inst_cellmath__24_0_I603 (.CO(N1494), .S(N1493), .A(N1488), .B(N1486), .CI(N1459));
ADDFX1 inst_cellmath__24_0_I604 (.CO(N1496), .S(N1495), .A(N1480), .B(N1456), .CI(N1477));
ADDFX1 arith_dfa_A_I2890 (.CO(N1499), .S(N6528), .A(N1493), .B(N1465), .CI(N1467));
ADDFX1 arith_dfa_A_I2891 (.CO(N1498), .S(N1497), .A(N1495), .B(N1472), .CI(N6528));
ADDHX1 inst_cellmath__24_0_I606 (.CO(N1501), .S(N1500), .A(N1094), .B(N427));
ADDFX1 arith_dfa_A_I2892 (.CO(N1504), .S(N6541), .A(N1476), .B(N487), .CI(N547));
ADDFX1 arith_dfa_A_I2893 (.CO(N1503), .S(N1502), .A(N1487), .B(N1479), .CI(N6541));
ADDFX1 arith_dfa_A_I2894 (.CO(N1507), .S(N6554), .A(N667), .B(N607), .CI(N727));
ADDFX1 arith_dfa_A_I2895 (.CO(N1506), .S(N1505), .A(N1489), .B(N1482), .CI(N6554));
ADDFX1 arith_dfa_A_I2896 (.CO(N1510), .S(N6567), .A(N847), .B(N787), .CI(N907));
ADDFX1 arith_dfa_A_I2897 (.CO(N1509), .S(N1508), .A(N967), .B(N1500), .CI(N6567));
ADDFX1 inst_cellmath__24_0_I610 (.CO(N1515), .S(N1514), .A(N1478), .B(N1027), .CI(N1481));
ADDFX1 inst_cellmath__24_0_I611 (.CO(N1517), .S(N1516), .A(N1508), .B(N1502), .CI(N1505));
ADDFX1 inst_cellmath__24_0_I612 (.CO(N1522), .S(N1521), .A(N1514), .B(N1494), .CI(N1496));
ADDFX1 inst_cellmath__24_0_I613 (.CO(N1524), .S(N1523), .A(N1499), .B(N1516), .CI(N1521));
ADDFX1 inst_cellmath__24_0_I614 (.CO(N1526), .S(N1525), .A(N1096), .B(N1093), .CI(N489));
ADDFX1 arith_dfa_A_I2898 (.CO(N1529), .S(N6580), .A(N429), .B(N549), .CI(N609));
ADDFX1 arith_dfa_A_I2899 (.CO(N1528), .S(N1527), .A(N1510), .B(N1507), .CI(N6580));
ADDFX1 arith_dfa_A_I2900 (.CO(N1532), .S(N6593), .A(N729), .B(N669), .CI(N789));
ADDFX1 arith_dfa_A_I2901 (.CO(N1531), .S(N1530), .A(N1501), .B(N1504), .CI(N6593));
ADDFX1 arith_dfa_A_I2902 (.CO(N1535), .S(N6606), .A(N909), .B(N849), .CI(N969));
ADDFX1 arith_dfa_A_I2903 (.CO(N1534), .S(N1533), .A(N1525), .B(N1029), .CI(N6606));
ADDFX1 arith_dfa_A_I2904 (.CO(N1538), .S(N6619), .A(N1506), .B(N1503), .CI(N1509));
ADDFX1 arith_dfa_A_I2905 (.CO(N1537), .S(N1536), .A(N1530), .B(N1515), .CI(N6619));
ADDFX1 inst_cellmath__24_0_I619 (.CO(N1543), .S(N1542), .A(N1533), .B(N1527), .CI(N1517));
ADDFX1 inst_cellmath__24_0_I620 (.CO(N1545), .S(N1544), .A(N1542), .B(N1522), .CI(N1536));
INVXL fap1_A_I2906 (.Y(N6636), .A(N1095));
ADDFX1 fap1_A_I2907 (.CO(N1547), .S(N1546), .A(N491), .B(N1098), .CI(N6636));
ADDFX1 arith_dfa_A_I2908 (.CO(N1552), .S(N6641), .A(N611), .B(N551), .CI(N671));
ADDFX1 arith_dfa_A_I2909 (.CO(N1551), .S(N1550), .A(N1535), .B(N1532), .CI(N6641));
ADDFX1 arith_dfa_A_I2910 (.CO(N1555), .S(N6654), .A(N791), .B(N731), .CI(N851));
ADDFX1 arith_dfa_A_I2911 (.CO(N1554), .S(N1553), .A(N1526), .B(N1529), .CI(N6654));
ADDFX1 inst_cellmath__24_0_I624 (.CO(N1560), .S(N1559), .A(N971), .B(N911), .CI(N1031));
ADDFX1 inst_cellmath__24_0_I625 (.CO(N1562), .S(N1561), .A(N1559), .B(N1212), .CI(N1546));
ADDFX1 arith_dfa_A_I2912 (.CO(N1565), .S(N6667), .A(N1531), .B(N1528), .CI(N1534));
ADDFX1 arith_dfa_A_I2913 (.CO(N1564), .S(N1563), .A(N1550), .B(N1538), .CI(N6667));
ADDFX1 inst_cellmath__24_0_I627 (.CO(N1570), .S(N1569), .A(N1553), .B(N1561), .CI(N1537));
ADDFX1 inst_cellmath__24_0_I628 (.CO(N1572), .S(N1571), .A(N1563), .B(N1543), .CI(N1569));
INVXL fap1_A_I2914 (.Y(N6684), .A(N1097));
ADDFX1 fap1_A_I2915 (.CO(N1574), .S(N1573), .A(N1100), .B(N1095), .CI(N6684));
ADDFX1 arith_dfa_A_I2916 (.CO(N1579), .S(N6689), .A(N493), .B(N553), .CI(N613));
ADDFX1 arith_dfa_A_I2917 (.CO(N1578), .S(N1577), .A(N1560), .B(N1547), .CI(N6689));
ADDFX1 arith_dfa_A_I2918 (.CO(N1582), .S(N6702), .A(N733), .B(N673), .CI(N793));
ADDFX1 arith_dfa_A_I2919 (.CO(N1581), .S(N1580), .A(N1555), .B(N1552), .CI(N6702));
ADDFX1 arith_dfa_A_I2920 (.CO(N1585), .S(N6715), .A(N913), .B(N853), .CI(N973));
ADDFX1 arith_dfa_A_I2921 (.CO(N1584), .S(N1583), .A(N1033), .B(N1573), .CI(N6715));
ADDFX1 arith_dfa_A_I2922 (.CO(N1588), .S(N6728), .A(N1562), .B(N1551), .CI(N1554));
ADDFX1 arith_dfa_A_I2923 (.CO(N1587), .S(N1586), .A(N1580), .B(N1565), .CI(N6728));
ADDFX1 inst_cellmath__24_0_I634 (.CO(N1593), .S(N1592), .A(N1583), .B(N1577), .CI(N1564));
ADDFX1 inst_cellmath__24_0_I635 (.CO(N1595), .S(N1594), .A(N1570), .B(N1586), .CI(N1592));
ADDFX1 inst_cellmath__24_0_I636 (.CO(N1597), .S(N1596), .A(N1097), .B(N1099), .CI(N1102));
ADDFX1 arith_dfa_A_I2924 (.CO(N1600), .S(N6741), .A(N615), .B(N555), .CI(N675));
ADDFX1 arith_dfa_A_I2925 (.CO(N1599), .S(N1598), .A(N1585), .B(N1582), .CI(N6741));
ADDFX1 arith_dfa_A_I2926 (.CO(N1603), .S(N6754), .A(N795), .B(N735), .CI(N855));
ADDFX1 arith_dfa_A_I2927 (.CO(N1602), .S(N1601), .A(N1574), .B(N1579), .CI(N6754));
ADDFX1 arith_dfa_A_I2928 (.CO(N1606), .S(N6767), .A(N975), .B(N915), .CI(N1035));
ADDFX1 arith_dfa_A_I2929 (.CO(N1605), .S(N1604), .A(N1213), .B(N1596), .CI(N6767));
ADDFX1 arith_dfa_A_I2930 (.CO(N1609), .S(N6780), .A(N1581), .B(N1578), .CI(N1584));
ADDFX1 arith_dfa_A_I2931 (.CO(N1608), .S(N1607), .A(N1598), .B(N1588), .CI(N6780));
ADDFX1 inst_cellmath__24_0_I641 (.CO(N1614), .S(N1613), .A(N1604), .B(N1601), .CI(N1587));
ADDFX1 inst_cellmath__24_0_I642 (.CO(N1616), .S(N1615), .A(N1593), .B(N1607), .CI(N1613));
INVXL fap1_A_I2932 (.Y(N6797), .A(N1101));
ADDFX1 fap1_A_I2933 (.CO(N1618), .S(N1617), .A(N617), .B(N1104), .CI(N6797));
ADDFX1 inst_cellmath__24_0_I644 (.CO(N1622), .S(N1621), .A(N737), .B(N677), .CI(N557));
ADDFX1 arith_dfa_A_I2934 (.CO(N1625), .S(N6802), .A(N857), .B(N797), .CI(N917));
ADDFX1 arith_dfa_A_I2935 (.CO(N1624), .S(N1623), .A(N1603), .B(N1600), .CI(N6802));
ADDFX1 arith_dfa_A_I2936 (.CO(N1628), .S(N6815), .A(N1037), .B(N977), .CI(N1597));
ADDFX1 arith_dfa_A_I2937 (.CO(N1627), .S(N1626), .A(N1621), .B(N1617), .CI(N6815));
ADDFX1 inst_cellmath__24_0_I647 (.CO(N1633), .S(N1632), .A(N1605), .B(N1606), .CI(N1599));
ADDFX1 inst_cellmath__24_0_I648 (.CO(N1635), .S(N1634), .A(N1623), .B(N1602), .CI(N1626));
ADDFX1 inst_cellmath__24_0_I649 (.CO(N1640), .S(N1639), .A(N1632), .B(N1609), .CI(N1634));
ADDFX1 inst_cellmath__24_0_I650 (.CO(N1642), .S(N1641), .A(N1614), .B(N1608), .CI(N1639));
ADDFX1 arith_dfa_A_I2938 (.CO(N1645), .S(N6828), .A(N1101), .B(N1103), .CI(N1106));
ADDFX1 arith_dfa_A_I2939 (.CO(N1644), .S(N1643), .A(N619), .B(N1214), .CI(N6828));
ADDFX1 arith_dfa_A_I2940 (.CO(N1648), .S(N6841), .A(N739), .B(N679), .CI(N799));
ADDFX1 arith_dfa_A_I2941 (.CO(N1647), .S(N1646), .A(N1622), .B(N1618), .CI(N6841));
ADDFX1 arith_dfa_A_I2942 (.CO(N1651), .S(N6854), .A(N919), .B(N859), .CI(N979));
ADDFX1 arith_dfa_A_I2943 (.CO(N1650), .S(N1649), .A(N1039), .B(N1625), .CI(N6854));
ADDFX1 inst_cellmath__24_0_I654 (.CO(N1656), .S(N1655), .A(N1643), .B(N1628), .CI(N1624));
ADDFX1 inst_cellmath__24_0_I655 (.CO(N1658), .S(N1657), .A(N1649), .B(N1627), .CI(N1646));
ADDFX1 arith_dfa_A_I2944 (.CO(N1661), .S(N6867), .A(N1655), .B(N1633), .CI(N1635));
ADDFX1 arith_dfa_A_I2945 (.CO(N1660), .S(N1659), .A(N1657), .B(N1640), .CI(N6867));
INVXL fap1_A_I2946 (.Y(N6884), .A(N1105));
ADDFX1 fap1_A_I2947 (.CO(N1663), .S(N1662), .A(N681), .B(N1108), .CI(N6884));
ADDFX1 arith_dfa_A_I2948 (.CO(N1668), .S(N6889), .A(N621), .B(N741), .CI(N801));
ADDFX1 arith_dfa_A_I2949 (.CO(N1667), .S(N1666), .A(N1651), .B(N1648), .CI(N6889));
ADDFX1 inst_cellmath__24_0_I659 (.CO(N1673), .S(N1672), .A(N921), .B(N861), .CI(N981));
ADDFX1 inst_cellmath__24_0_I660 (.CO(N1675), .S(N1674), .A(N1645), .B(N1041), .CI(N1672));
ADDFX1 inst_cellmath__24_0_I661 (.CO(N1680), .S(N1679), .A(N1644), .B(N1662), .CI(N1650));
ADDFX1 inst_cellmath__24_0_I662 (.CO(N1682), .S(N1681), .A(N1674), .B(N1647), .CI(N1666));
ADDFX1 inst_cellmath__24_0_I663 (.CO(N1687), .S(N1686), .A(N1679), .B(N1656), .CI(N1658));
ADDFX1 inst_cellmath__24_0_I664 (.CO(N1689), .S(N1688), .A(N1661), .B(N1681), .CI(N1686));
ADDFX1 inst_cellmath__24_0_I665 (.CO(N1691), .S(N1690), .A(N1105), .B(N1107), .CI(N1110));
ADDFX1 arith_dfa_A_I2950 (.CO(N1694), .S(N6902), .A(N743), .B(N683), .CI(N803));
ADDFX1 arith_dfa_A_I2951 (.CO(N1693), .S(N1692), .A(N1673), .B(N1663), .CI(N6902));
ADDFX1 arith_dfa_A_I2952 (.CO(N1697), .S(N6915), .A(N923), .B(N863), .CI(N983));
ADDFX1 arith_dfa_A_I2953 (.CO(N1696), .S(N1695), .A(N1690), .B(N1668), .CI(N6915));
ADDFX1 inst_cellmath__24_0_I668 (.CO(N1702), .S(N1701), .A(N1215), .B(N1043), .CI(N1667));
ADDFX1 inst_cellmath__24_0_I669 (.CO(N1704), .S(N1703), .A(N1695), .B(N1675), .CI(N1692));
ADDFX1 arith_dfa_A_I2954 (.CO(N1707), .S(N6928), .A(N1701), .B(N1680), .CI(N1682));
ADDFX1 arith_dfa_A_I2955 (.CO(N1706), .S(N1705), .A(N1703), .B(N1687), .CI(N6928));
INVXL fap1_A_I2956 (.Y(N6945), .A(N1109));
ADDFX1 fap1_A_I2957 (.CO(N1709), .S(N1708), .A(N745), .B(N1112), .CI(N6945));
ADDFX1 inst_cellmath__24_0_I672 (.CO(N1713), .S(N1712), .A(N865), .B(N805), .CI(N685));
ADDFX1 arith_dfa_A_I2958 (.CO(N1716), .S(N6950), .A(N985), .B(N925), .CI(N1045));
ADDFX1 arith_dfa_A_I2959 (.CO(N1715), .S(N1714), .A(N1697), .B(N1694), .CI(N6950));
ADDFX1 inst_cellmath__24_0_I674 (.CO(N1721), .S(N1720), .A(N1712), .B(N1691), .CI(N1708));
ADDFX1 inst_cellmath__24_0_I675 (.CO(N1723), .S(N1722), .A(N1696), .B(N1693), .CI(N1720));
ADDFX1 inst_cellmath__24_0_I676 (.CO(N1728), .S(N1727), .A(N1702), .B(N1714), .CI(N1704));
ADDFX1 inst_cellmath__24_0_I677 (.CO(N1730), .S(N1729), .A(N1707), .B(N1722), .CI(N1727));
ADDFX1 arith_dfa_A_I2960 (.CO(N1733), .S(N6963), .A(N1109), .B(N1111), .CI(N1114));
ADDFX1 arith_dfa_A_I2961 (.CO(N1732), .S(N1731), .A(N747), .B(N1216), .CI(N6963));
ADDFX1 arith_dfa_A_I2962 (.CO(N1736), .S(N6976), .A(N867), .B(N807), .CI(N927));
ADDFX1 arith_dfa_A_I2963 (.CO(N1735), .S(N1734), .A(N1713), .B(N1709), .CI(N6976));
ADDFX1 inst_cellmath__24_0_I680 (.CO(N1741), .S(N1740), .A(N1047), .B(N987), .CI(N1716));
ADDFX1 inst_cellmath__24_0_I681 (.CO(N1743), .S(N1742), .A(N1740), .B(N1731), .CI(N1715));
ADDFX1 inst_cellmath__24_0_I682 (.CO(N1748), .S(N1747), .A(N1734), .B(N1721), .CI(N1742));
ADDFX1 inst_cellmath__24_0_I683 (.CO(N1750), .S(N1749), .A(N1728), .B(N1723), .CI(N1747));
INVXL fap1_A_I2964 (.Y(N6993), .A(N1113));
ADDFX1 fap1_A_I2965 (.CO(N1752), .S(N1751), .A(N809), .B(N1116), .CI(N6993));
ADDFX1 arith_dfa_A_I2966 (.CO(N1757), .S(N6998), .A(N749), .B(N869), .CI(N929));
ADDFX1 arith_dfa_A_I2967 (.CO(N1756), .S(N1755), .A(N1733), .B(N1736), .CI(N6998));
ADDFX1 inst_cellmath__24_0_I686 (.CO(N1762), .S(N1761), .A(N1049), .B(N989), .CI(N1751));
ADDFX1 inst_cellmath__24_0_I687 (.CO(N1764), .S(N1763), .A(N1741), .B(N1732), .CI(N1735));
ADDFX1 arith_dfa_A_I2968 (.CO(N1767), .S(N7011), .A(N1755), .B(N1761), .CI(N1743));
ADDFX1 arith_dfa_A_I2969 (.CO(N1766), .S(N1765), .A(N1763), .B(N1748), .CI(N7011));
ADDFX1 inst_cellmath__24_0_I689 (.CO(N1769), .S(N1768), .A(N1113), .B(N1115), .CI(N1118));
ADDFX1 arith_dfa_A_I2970 (.CO(N1772), .S(N7024), .A(N871), .B(N811), .CI(N931));
ADDFX1 arith_dfa_A_I2971 (.CO(N1771), .S(N1770), .A(N1757), .B(N1752), .CI(N7024));
ADDFX1 inst_cellmath__24_0_I691 (.CO(N1777), .S(N1776), .A(N1051), .B(N991), .CI(N1217));
ADDFX1 inst_cellmath__24_0_I692 (.CO(N1779), .S(N1778), .A(N1776), .B(N1768), .CI(N1756));
ADDFX1 inst_cellmath__24_0_I693 (.CO(N1784), .S(N1783), .A(N1770), .B(N1762), .CI(N1764));
ADDFX1 inst_cellmath__24_0_I694 (.CO(N1786), .S(N1785), .A(N1767), .B(N1778), .CI(N1783));
INVXL fap1_A_I2972 (.Y(N7041), .A(N1117));
ADDFX1 fap1_A_I2973 (.CO(N1788), .S(N1787), .A(N873), .B(N1120), .CI(N7041));
ADDFX1 inst_cellmath__24_0_I696 (.CO(N1792), .S(N1791), .A(N993), .B(N933), .CI(N813));
ADDFX1 inst_cellmath__24_0_I697 (.CO(N1797), .S(N1796), .A(N1769), .B(N1053), .CI(N1772));
ADDFX1 inst_cellmath__24_0_I698 (.CO(N1799), .S(N1798), .A(N1791), .B(N1777), .CI(N1787));
ADDFX1 arith_dfa_A_I2974 (.CO(N1802), .S(N7046), .A(N1771), .B(N1796), .CI(N1798));
ADDFX1 arith_dfa_A_I2975 (.CO(N1801), .S(N1800), .A(N1779), .B(N1784), .CI(N7046));
ADDFX1 arith_dfa_A_I2976 (.CO(N1805), .S(N7059), .A(N1117), .B(N1119), .CI(N1122));
ADDFX1 arith_dfa_A_I2977 (.CO(N1804), .S(N1803), .A(N875), .B(N1218), .CI(N7059));
ADDFX1 arith_dfa_A_I2978 (.CO(N1808), .S(N7072), .A(N995), .B(N935), .CI(N1055));
ADDFX1 arith_dfa_A_I2979 (.CO(N1807), .S(N1806), .A(N1792), .B(N1788), .CI(N7072));
ADDFX1 arith_dfa_A_I2980 (.CO(N1811), .S(N7085), .A(N1803), .B(N1797), .CI(N1799));
ADDFX1 arith_dfa_A_I2981 (.CO(N1810), .S(N1809), .A(N1806), .B(N1802), .CI(N7085));
INVXL fap1_A_I2982 (.Y(N7102), .A(N1121));
ADDFX1 fap1_A_I2983 (.CO(N1813), .S(N1812), .A(N937), .B(N1124), .CI(N7102));
ADDFX1 arith_dfa_A_I2984 (.CO(N1818), .S(N7107), .A(N877), .B(N997), .CI(N1057));
ADDFX1 arith_dfa_A_I2985 (.CO(N1817), .S(N1816), .A(N1805), .B(N1808), .CI(N7107));
ADDFX1 inst_cellmath__24_0_I705 (.CO(N1823), .S(N1822), .A(N1804), .B(N1812), .CI(N1807));
ADDFX1 inst_cellmath__24_0_I706 (.CO(N1825), .S(N1824), .A(N1811), .B(N1816), .CI(N1822));
ADDFX1 inst_cellmath__24_0_I707 (.CO(N1827), .S(N1826), .A(N1121), .B(N1123), .CI(N1126));
ADDFX1 arith_dfa_A_I2986 (.CO(N1830), .S(N7120), .A(N999), .B(N939), .CI(N1059));
ADDFX1 arith_dfa_A_I2987 (.CO(N1829), .S(N1828), .A(N1818), .B(N1813), .CI(N7120));
ADDFX1 inst_cellmath__24_0_I709 (.CO(N1835), .S(N1834), .A(N1826), .B(N1219), .CI(N1817));
ADDFX1 inst_cellmath__24_0_I710 (.CO(N1837), .S(N1836), .A(N1823), .B(N1828), .CI(N1834));
INVXL fap1_A_I2988 (.Y(N7137), .A(N1125));
ADDFX1 fap1_A_I2989 (.CO(N1839), .S(N1838), .A(N1001), .B(N1128), .CI(N7137));
ADDFX1 inst_cellmath__24_0_I712 (.CO(N1843), .S(N1842), .A(N941), .B(N1061), .CI(N1827));
ADDFX1 arith_dfa_A_I2990 (.CO(N1846), .S(N7142), .A(N1838), .B(N1830), .CI(N1842));
ADDFX1 arith_dfa_A_I2991 (.CO(N1845), .S(N1844), .A(N1835), .B(N1829), .CI(N7142));
ADDFX1 arith_dfa_A_I2992 (.CO(N1849), .S(N7155), .A(N1125), .B(N1127), .CI(N1130));
ADDFX1 arith_dfa_A_I2993 (.CO(N1848), .S(N1847), .A(N1003), .B(N1220), .CI(N7155));
ADDFX1 inst_cellmath__24_0_I715 (.CO(N1854), .S(N1853), .A(N1839), .B(N1063), .CI(N1843));
ADDFX1 inst_cellmath__24_0_I716 (.CO(N1856), .S(N1855), .A(N1853), .B(N1847), .CI(N1846));
INVXL fap1_A_I2994 (.Y(N7172), .A(N1129));
ADDFX1 fap1_A_I2995 (.CO(N1858), .S(N1857), .A(N1065), .B(N1132), .CI(N7172));
ADDFX1 inst_cellmath__24_0_I718 (.CO(N1865), .S(N1864), .A(N1849), .B(N1005), .CI(N1857));
ADDFX1 inst_cellmath__24_0_I719 (.CO(N1867), .S(N1866), .A(N1854), .B(N1848), .CI(N1864));
ADDFX1 inst_cellmath__24_0_I720 (.CO(N1869), .S(N1868), .A(N1129), .B(N1131), .CI(N1134));
ADDFX1 inst_cellmath__24_0_I721 (.CO(N1874), .S(N1873), .A(N1221), .B(N1067), .CI(N1868));
ADDFX1 inst_cellmath__24_0_I722 (.CO(N1876), .S(N1875), .A(N1873), .B(N1858), .CI(N1865));
INVXL fap1_A_I2996 (.Y(N7181), .A(N1133));
ADDFX1 fap1_A_I2997 (.CO(N1878), .S(N1877), .A(N1069), .B(N1136), .CI(N7181));
ADDFX1 inst_cellmath__24_0_I724 (.CO(N1882), .S(N1881), .A(N1877), .B(N1869), .CI(N1874));
ADDFX1 inst_cellmath__24_0_I725 (.CO(N1887), .S(N1886), .A(N1133), .B(N1135), .CI(N1138));
ADDFX1 inst_cellmath__24_0_I726 (.CO(N1889), .S(N1888), .A(N1886), .B(N1222), .CI(N1878));
ADDFX1 inst_cellmath__24_0_I728 (.CO(N1895), .S(N1894), .A(N7692), .B(N1140), .CI(N1887));
XNOR2X1 inst_cellmath__24_0_I730 (.Y(N1900), .A(N1144), .B(N7692));
AND2XL inst_cellmath__24_0_I731 (.Y(N1902), .A(inst_cellmath__24_0_in0[1]), .B(N381));
NOR2XL inst_cellmath__24_0_I733 (.Y(N1904), .A(N445), .B(N1223));
NAND2XL inst_cellmath__24_0_I734 (.Y(N1905), .A(N445), .B(N1223));
NOR2XL inst_cellmath__24_0_I735 (.Y(N1906), .A(N1224), .B(N1225));
NAND2XL inst_cellmath__24_0_I736 (.Y(N1907), .A(N1224), .B(N1225));
NOR2XL inst_cellmath__24_0_I737 (.Y(N1908), .A(N1227), .B(N1229));
NAND2XL inst_cellmath__24_0_I738 (.Y(N1909), .A(N1227), .B(N1229));
NOR2XL inst_cellmath__24_0_I739 (.Y(N1910), .A(N1230), .B(N1233));
NAND2XL inst_cellmath__24_0_I740 (.Y(N1911), .A(N1230), .B(N1233));
NOR2XL inst_cellmath__24_0_I741 (.Y(N1912), .A(N1234), .B(N1237));
NAND2XL inst_cellmath__24_0_I742 (.Y(N1913), .A(N1234), .B(N1237));
NOR2XL inst_cellmath__24_0_I743 (.Y(N1914), .A(N1238), .B(N1247));
NAND2XL inst_cellmath__24_0_I744 (.Y(N1915), .A(N1238), .B(N1247));
NOR2XL inst_cellmath__24_0_I745 (.Y(N1916), .A(N1248), .B(N1253));
NAND2XL inst_cellmath__24_0_I746 (.Y(N1917), .A(N1248), .B(N1253));
NOR2XL inst_cellmath__24_0_I747 (.Y(N1918), .A(N1254), .B(N1265));
NAND2XL inst_cellmath__24_0_I748 (.Y(N1919), .A(N1254), .B(N1265));
NOR2XL inst_cellmath__24_0_I749 (.Y(N1920), .A(N1266), .B(N1277));
NAND2XL inst_cellmath__24_0_I750 (.Y(N1921), .A(N1266), .B(N1277));
NOR2XL inst_cellmath__24_0_I751 (.Y(N1922), .A(N1278), .B(N1289));
NAND2XL inst_cellmath__24_0_I752 (.Y(N1923), .A(N1278), .B(N1289));
NOR2XL inst_cellmath__24_0_I753 (.Y(N1924), .A(N1290), .B(N1303));
NAND2XL inst_cellmath__24_0_I754 (.Y(N1925), .A(N1290), .B(N1303));
NOR2XL inst_cellmath__24_0_I755 (.Y(N1926), .A(N1304), .B(N1321));
NAND2XL inst_cellmath__24_0_I756 (.Y(N1927), .A(N1304), .B(N1321));
NOR2XL inst_cellmath__24_0_I757 (.Y(N1928), .A(N1322), .B(N1336));
NAND2XL inst_cellmath__24_0_I758 (.Y(N1929), .A(N1322), .B(N1336));
NOR2XL inst_cellmath__24_0_I759 (.Y(N1930), .A(N1337), .B(N1351));
NAND2XL inst_cellmath__24_0_I760 (.Y(N1931), .A(N1337), .B(N1351));
NOR2X1 inst_cellmath__24_0_I761 (.Y(N1932), .A(N1352), .B(N1372));
NAND2XL inst_cellmath__24_0_I762 (.Y(N1933), .A(N1352), .B(N1372));
NOR2XL inst_cellmath__24_0_I763 (.Y(N1934), .A(N1373), .B(N1393));
NAND2X1 inst_cellmath__24_0_I764 (.Y(N1935), .A(N1373), .B(N1393));
NOR2XL inst_cellmath__24_0_I765 (.Y(N1936), .A(N1394), .B(N1410));
NAND2XL inst_cellmath__24_0_I766 (.Y(N1937), .A(N1394), .B(N1410));
AND2XL inst_cellmath__24_0_I769 (.Y(N1940), .A(N1903), .B(N1902));
INVXL inst_cellmath__24_0_I3408 (.Y(N7910), .A(N1904));
INVXL inst_cellmath__24_0_I3409 (.Y(N7911), .A(N1905));
OAI21XL inst_cellmath__24_0_I777 (.Y(N1950), .A0(N7911), .A1(N1940), .B0(N7910));
AOI21XL inst_cellmath__24_0_I785 (.Y(N1958), .A0(N1907), .A1(N1950), .B0(N1906));
INVXL inst_cellmath__24_0_I3415 (.Y(N7917), .A(N1908));
INVXL inst_cellmath__24_0_I3416 (.Y(N7918), .A(N1909));
OAI21XL inst_cellmath__24_0_I797 (.Y(N1970), .A0(N7918), .A1(N1958), .B0(N7917));
AOI21XL inst_cellmath__24_0_I809 (.Y(N1982), .A0(N1911), .A1(N1970), .B0(N1910));
INVXL inst_cellmath__24_0_I3426 (.Y(N7928), .A(N1912));
INVXL inst_cellmath__24_0_I3427 (.Y(N7929), .A(N1913));
OAI21X1 inst_cellmath__24_0_I825 (.Y(N1998), .A0(N7929), .A1(N1982), .B0(N7928));
AO21XL inst_cellmath__24_0_I3535 (.Y(N7940), .A0(N1917), .A1(N1914), .B0(N1916));
AOI21XL inst_cellmath__24_0_I849 (.Y(N2022), .A0(N1915), .A1(N1998), .B0(N1914));
AOI31X1 inst_cellmath__24_0_I3557 (.Y(N2024), .A0(N1917), .A1(N1915), .A2(N1998), .B0(N7940));
INVXL inst_cellmath__24_0_I3447 (.Y(N7949), .A(N1918));
INVXL inst_cellmath__24_0_I3448 (.Y(N7950), .A(N1919));
OAI21X1 inst_cellmath__24_0_I873 (.Y(N2046), .A0(N7950), .A1(N2024), .B0(N7949));
AO21XL inst_cellmath__24_0_I3538 (.Y(N7964), .A0(N1923), .A1(N1920), .B0(N1922));
AND2XL inst_cellmath__24_0_I3539 (.Y(N7965), .A(N1923), .B(N1921));
AOI21XL inst_cellmath__24_0_I903 (.Y(N2076), .A0(N1921), .A1(N2046), .B0(N1920));
AOI21X1 inst_cellmath__24_0_I905 (.Y(N2078), .A0(N7965), .A1(N2046), .B0(N7964));
INVXL inst_cellmath__24_0_I3475 (.Y(N7977), .A(N1925));
AOI21XL inst_cellmath__24_0_I909 (.Y(N2082), .A0(N1927), .A1(N1924), .B0(N1926));
NAND2XL inst_cellmath__24_0_I910 (.Y(N2083), .A(N1927), .B(N1925));
OAI21X2 inst_cellmath__24_0_I937 (.Y(N2110), .A0(N2083), .A1(N2078), .B0(N2082));
AO21XL inst_cellmath__24_0_I3541 (.Y(N7994), .A0(N1931), .A1(N1928), .B0(N1930));
AND2XL inst_cellmath__24_0_I3542 (.Y(N7995), .A(N1931), .B(N1929));
NOR2XL andori2bb1_A_I3579 (.Y(N8028), .A(N7977), .B(N2078));
NOR2XL andori2bb1_A_I3580 (.Y(N8008), .A(N8028), .B(N1924));
AOI21XL inst_cellmath__24_0_I975 (.Y(N2148), .A0(N1929), .A1(N2110), .B0(N1928));
AOI21X2 inst_cellmath__24_0_I977 (.Y(N2150), .A0(N7995), .A1(N2110), .B0(N7994));
AOI21XL inst_cellmath__24_0_I981 (.Y(N2154), .A0(N1935), .A1(N1932), .B0(N1934));
NAND2XL inst_cellmath__24_0_I982 (.Y(N2155), .A(N1935), .B(N1933));
INVXL inst_cellmath__24_0_I3511 (.Y(N8013), .A(N1937));
INVXL inst_cellmath__24_0_I3516 (.Y(N8018), .A(N1932));
INVXL inst_cellmath__24_0_I3517 (.Y(N8019), .A(N1933));
NOR2XL andori2bb1_A_I3581 (.Y(N8035), .A(N8013), .B(N2154));
NOR2XL andori2bb1_A_I3582 (.Y(N8022), .A(N8035), .B(N1936));
OAI21XL inst_cellmath__24_0_I1029 (.Y(N2202), .A0(N8019), .A1(N2150), .B0(N8018));
OAI21XL inst_cellmath__24_0_I1031 (.Y(N2204), .A0(N2155), .A1(N2150), .B0(N2154));
OAI31X1 inst_cellmath__24_0_I3573 (.Y(N2287), .A0(N8013), .A1(N2155), .A2(N2150), .B0(N8022));
NAND2BXL inst_cellmath__24_0_I1043 (.Y(N2218), .AN(N1904), .B(N1905));
NAND2BXL inst_cellmath__24_0_I1046 (.Y(N2221), .AN(N1906), .B(N1907));
NAND2BXL inst_cellmath__24_0_I1049 (.Y(N2224), .AN(N1908), .B(N1909));
NAND2BXL inst_cellmath__24_0_I1052 (.Y(N2227), .AN(N1910), .B(N1911));
NAND2BXL inst_cellmath__24_0_I1055 (.Y(N2230), .AN(N1912), .B(N1913));
NAND2BXL inst_cellmath__24_0_I1058 (.Y(N2233), .AN(N1914), .B(N1915));
NAND2BXL inst_cellmath__24_0_I1061 (.Y(N2236), .AN(N1916), .B(N1917));
NAND2BXL inst_cellmath__24_0_I1064 (.Y(N2239), .AN(N1918), .B(N1919));
NAND2BXL inst_cellmath__24_0_I1067 (.Y(N2242), .AN(N1920), .B(N1921));
NAND2BXL inst_cellmath__24_0_I1070 (.Y(N2245), .AN(N1922), .B(N1923));
NAND2BXL inst_cellmath__24_0_I1073 (.Y(N2248), .AN(N1924), .B(N1925));
NAND2BXL inst_cellmath__24_0_I1076 (.Y(N2251), .AN(N1926), .B(N1927));
NAND2BXL inst_cellmath__24_0_I1079 (.Y(N2254), .AN(N1928), .B(N1929));
NAND2BXL inst_cellmath__24_0_I1082 (.Y(N2257), .AN(N1930), .B(N1931));
NAND2BXL inst_cellmath__24_0_I1085 (.Y(N2260), .AN(N1932), .B(N1933));
NAND2BXL inst_cellmath__24_0_I1088 (.Y(N2263), .AN(N1934), .B(N1935));
NAND2BXL inst_cellmath__24_0_I1091 (.Y(N2266), .AN(N1936), .B(N1937));
XOR2XL inst_cellmath__24_0_I1092 (.Y(inst_cellmath__24_0_out0[0]), .A(inst_cellmath__24_0_in0[1]), .B(N381));
XOR2XL inst_cellmath__24_0_I3547 (.Y(inst_cellmath__24_0_out0[1]), .A(N1902), .B(N1903));
XNOR2X1 inst_cellmath__24_0_I1094 (.Y(inst_cellmath__24_0_out0[2]), .A(N1940), .B(N2218));
XOR2XL inst_cellmath__24_0_I3548 (.Y(inst_cellmath__24_0_out0[3]), .A(N1950), .B(N2221));
XNOR2X1 inst_cellmath__24_0_I1096 (.Y(inst_cellmath__24_0_out0[4]), .A(N1958), .B(N2224));
XOR2XL inst_cellmath__24_0_I3549 (.Y(inst_cellmath__24_0_out0[5]), .A(N1970), .B(N2227));
XNOR2X1 inst_cellmath__24_0_I1098 (.Y(inst_cellmath__24_0_out0[6]), .A(N1982), .B(N2230));
XOR2XL inst_cellmath__24_0_I3550 (.Y(inst_cellmath__24_0_out0[7]), .A(N1998), .B(N2233));
XNOR2X1 inst_cellmath__24_0_I1100 (.Y(inst_cellmath__24_0_out0[8]), .A(N2022), .B(N2236));
XNOR2X1 inst_cellmath__24_0_I1101 (.Y(inst_cellmath__24_0_out0[9]), .A(N2024), .B(N2239));
XOR2XL inst_cellmath__24_0_I3551 (.Y(inst_cellmath__24_0_out0[10]), .A(N2046), .B(N2242));
XNOR2X1 inst_cellmath__24_0_I1103 (.Y(inst_cellmath__24_0_out0[11]), .A(N2076), .B(N2245));
XNOR2X1 inst_cellmath__24_0_I1104 (.Y(inst_cellmath__24_0_out0[12]), .A(N2078), .B(N2248));
XNOR2X1 inst_cellmath__24_0_I1105 (.Y(inst_cellmath__24_0_out0[13]), .A(N8008), .B(N2251));
XOR2XL inst_cellmath__24_0_I3552 (.Y(inst_cellmath__24_0_out0[14]), .A(N2110), .B(N2254));
XNOR2X1 inst_cellmath__24_0_I1107 (.Y(inst_cellmath__24_0_out0[15]), .A(N2148), .B(N2257));
XNOR2X1 inst_cellmath__24_0_I1108 (.Y(inst_cellmath__24_0_out0[16]), .A(N2150), .B(N2260));
XOR2XL inst_cellmath__24_0_I1109 (.Y(inst_cellmath__24_0_out0[17]), .A(N2202), .B(N2263));
XOR2XL inst_cellmath__24_0_I1110 (.Y(inst_cellmath__24_0_out0[18]), .A(N2204), .B(N2266));
OR2XL inst_cellmath__24_0_I1113 (.Y(N7186), .A(N1411), .B(N1428));
XOR2XL inst_cellmath__24_0_I1114 (.Y(N2290), .A(N1411), .B(N1428));
OR2XL inst_cellmath__24_0_I1115 (.Y(N7193), .A(N1429), .B(N1448));
XOR2XL inst_cellmath__24_0_I1116 (.Y(N2292), .A(N1429), .B(N1448));
XOR2XL inst_cellmath__24_0_I1118 (.Y(N2294), .A(N1449), .B(N1473));
XOR2XL inst_cellmath__24_0_I1120 (.Y(N2296), .A(N1474), .B(N1497));
OR2XL inst_cellmath__24_0_I1121 (.Y(N7214), .A(N1498), .B(N1523));
XOR2XL inst_cellmath__24_0_I1122 (.Y(N2298), .A(N1498), .B(N1523));
OR2XL inst_cellmath__24_0_I1123 (.Y(N7221), .A(N1524), .B(N1544));
XOR2XL inst_cellmath__24_0_I1124 (.Y(N2300), .A(N1524), .B(N1544));
OR2XL inst_cellmath__24_0_I1125 (.Y(N7228), .A(N1545), .B(N1571));
XOR2XL inst_cellmath__24_0_I1126 (.Y(N2302), .A(N1545), .B(N1571));
OR2XL inst_cellmath__24_0_I1127 (.Y(N7235), .A(N1572), .B(N1594));
XOR2XL inst_cellmath__24_0_I1128 (.Y(N2304), .A(N1572), .B(N1594));
OR2XL inst_cellmath__24_0_I1129 (.Y(N7242), .A(N1595), .B(N1615));
XOR2XL inst_cellmath__24_0_I1130 (.Y(N2306), .A(N1595), .B(N1615));
OR2XL inst_cellmath__24_0_I1131 (.Y(N7249), .A(N1616), .B(N1641));
XOR2XL inst_cellmath__24_0_I1132 (.Y(N2308), .A(N1616), .B(N1641));
OR2XL inst_cellmath__24_0_I1133 (.Y(N7256), .A(N1642), .B(N1659));
XOR2XL inst_cellmath__24_0_I1134 (.Y(N2310), .A(N1642), .B(N1659));
OR2XL inst_cellmath__24_0_I1135 (.Y(N7263), .A(N1660), .B(N1688));
XOR2XL inst_cellmath__24_0_I1136 (.Y(N2312), .A(N1660), .B(N1688));
OR2XL inst_cellmath__24_0_I1137 (.Y(N7270), .A(N1689), .B(N1705));
XOR2XL inst_cellmath__24_0_I1138 (.Y(N2314), .A(N1689), .B(N1705));
OR2XL inst_cellmath__24_0_I1139 (.Y(N7277), .A(N1706), .B(N1729));
XOR2XL inst_cellmath__24_0_I1140 (.Y(N2316), .A(N1706), .B(N1729));
OR2XL inst_cellmath__24_0_I1141 (.Y(N7284), .A(N1730), .B(N1749));
XOR2XL inst_cellmath__24_0_I1142 (.Y(N2318), .A(N1730), .B(N1749));
OR2XL inst_cellmath__24_0_I1143 (.Y(N7291), .A(N1750), .B(N1765));
XOR2XL inst_cellmath__24_0_I1144 (.Y(N2320), .A(N1750), .B(N1765));
OR2XL inst_cellmath__24_0_I1145 (.Y(N7298), .A(N1766), .B(N1785));
XOR2XL inst_cellmath__24_0_I1146 (.Y(N2322), .A(N1766), .B(N1785));
OR2XL inst_cellmath__24_0_I1147 (.Y(N7305), .A(N1786), .B(N1800));
XOR2XL inst_cellmath__24_0_I1148 (.Y(N2324), .A(N1786), .B(N1800));
OR2XL inst_cellmath__24_0_I1149 (.Y(N7312), .A(N1801), .B(N1809));
XOR2XL inst_cellmath__24_0_I1150 (.Y(N2326), .A(N1801), .B(N1809));
OR2XL inst_cellmath__24_0_I1151 (.Y(N7319), .A(N1810), .B(N1824));
XOR2XL inst_cellmath__24_0_I1152 (.Y(N2328), .A(N1810), .B(N1824));
OR2XL inst_cellmath__24_0_I1153 (.Y(N7326), .A(N1825), .B(N1836));
XOR2XL inst_cellmath__24_0_I1154 (.Y(N2330), .A(N1825), .B(N1836));
OR2XL inst_cellmath__24_0_I1155 (.Y(N7333), .A(N1837), .B(N1844));
XOR2XL inst_cellmath__24_0_I1156 (.Y(N2332), .A(N1837), .B(N1844));
OR2XL inst_cellmath__24_0_I1157 (.Y(N7340), .A(N1855), .B(N1845));
XOR2XL inst_cellmath__24_0_I1158 (.Y(N2334), .A(N1855), .B(N1845));
OR2XL inst_cellmath__24_0_I1159 (.Y(N7347), .A(N1856), .B(N1866));
XOR2XL inst_cellmath__24_0_I1160 (.Y(N2336), .A(N1856), .B(N1866));
OR2XL inst_cellmath__24_0_I1161 (.Y(N7354), .A(N1867), .B(N1875));
XOR2XL inst_cellmath__24_0_I1162 (.Y(N2338), .A(N1867), .B(N1875));
OR2XL inst_cellmath__24_0_I1163 (.Y(N7361), .A(N1881), .B(N1876));
XOR2XL inst_cellmath__24_0_I1164 (.Y(N2340), .A(N1881), .B(N1876));
OR2XL inst_cellmath__24_0_I1165 (.Y(N7368), .A(N1888), .B(N1882));
XOR2XL inst_cellmath__24_0_I1166 (.Y(N2342), .A(N1888), .B(N1882));
OR2XL inst_cellmath__24_0_I1167 (.Y(N7375), .A(N1894), .B(N1889));
XOR2XL inst_cellmath__24_0_I1168 (.Y(N2344), .A(N1894), .B(N1889));
XNOR2X1 inst_cellmath__24_0_I1170 (.Y(N2346), .A(N1895), .B(N1900));
OAI2BB1X1 inst_cellmath__24_0_I2999 (.Y(N2349), .A0N(N2290), .A1N(N2287), .B0(N7186));
OAI2BB1X1 inst_cellmath__24_0_I3001 (.Y(N2355), .A0N(N2292), .A1N(N2349), .B0(N7193));
OAI2BB2XL inst_cellmath__24_0_I3553 (.Y(N2363), .A0N(N2294), .A1N(N2355), .B0(N1449), .B1(N1473));
OAI2BB2XL inst_cellmath__24_0_I3554 (.Y(N2373), .A0N(N2296), .A1N(N2363), .B0(N1474), .B1(N1497));
OAI2BB1X1 inst_cellmath__24_0_I3007 (.Y(N2385), .A0N(N2298), .A1N(N2373), .B0(N7214));
OAI2BB1X1 inst_cellmath__24_0_I3009 (.Y(N2399), .A0N(N2300), .A1N(N2385), .B0(N7221));
OAI2BB1X1 inst_cellmath__24_0_I3011 (.Y(N2415), .A0N(N2302), .A1N(N2399), .B0(N7228));
OAI2BB1X1 inst_cellmath__24_0_I3013 (.Y(N2433), .A0N(N2304), .A1N(N2415), .B0(N7235));
OAI2BB1X1 inst_cellmath__24_0_I3015 (.Y(N2453), .A0N(N2306), .A1N(N2433), .B0(N7242));
OAI2BB1X1 inst_cellmath__24_0_I3017 (.Y(N2475), .A0N(N2308), .A1N(N2453), .B0(N7249));
OAI2BB1X1 inst_cellmath__24_0_I3019 (.Y(N2499), .A0N(N2310), .A1N(N2475), .B0(N7256));
OAI2BB1X1 inst_cellmath__24_0_I3021 (.Y(N2525), .A0N(N2312), .A1N(N2499), .B0(N7263));
OAI2BB1X1 inst_cellmath__24_0_I3023 (.Y(N2553), .A0N(N2314), .A1N(N2525), .B0(N7270));
OAI2BB1X1 inst_cellmath__24_0_I3025 (.Y(N2583), .A0N(N2316), .A1N(N2553), .B0(N7277));
OAI2BB1X1 inst_cellmath__24_0_I3027 (.Y(N2615), .A0N(N2318), .A1N(N2583), .B0(N7284));
OAI2BB1X1 inst_cellmath__24_0_I3029 (.Y(N2649), .A0N(N2320), .A1N(N2615), .B0(N7291));
OAI2BB1X1 inst_cellmath__24_0_I3031 (.Y(N2685), .A0N(N2322), .A1N(N2649), .B0(N7298));
OAI2BB1X1 inst_cellmath__24_0_I3033 (.Y(N2723), .A0N(N2324), .A1N(N2685), .B0(N7305));
OAI2BB1X1 inst_cellmath__24_0_I3035 (.Y(N2763), .A0N(N2326), .A1N(N2723), .B0(N7312));
OAI2BB1X1 inst_cellmath__24_0_I3037 (.Y(N2805), .A0N(N2328), .A1N(N2763), .B0(N7319));
OAI2BB1X1 inst_cellmath__24_0_I3039 (.Y(N2849), .A0N(N2330), .A1N(N2805), .B0(N7326));
OAI2BB1X1 inst_cellmath__24_0_I3041 (.Y(N2895), .A0N(N2332), .A1N(N2849), .B0(N7333));
OAI2BB1X1 inst_cellmath__24_0_I3043 (.Y(N2943), .A0N(N2334), .A1N(N2895), .B0(N7340));
OAI2BB1X1 inst_cellmath__24_0_I3045 (.Y(N2993), .A0N(N2336), .A1N(N2943), .B0(N7347));
OAI2BB1X1 inst_cellmath__24_0_I3047 (.Y(N3045), .A0N(N2338), .A1N(N2993), .B0(N7354));
OAI2BB1X1 inst_cellmath__24_0_I3049 (.Y(N3099), .A0N(N2340), .A1N(N3045), .B0(N7361));
OAI2BB1X1 inst_cellmath__24_0_I3051 (.Y(N3155), .A0N(N2342), .A1N(N3099), .B0(N7368));
OAI2BB1X1 inst_cellmath__24_0_I3053 (.Y(N3213), .A0N(N2344), .A1N(N3155), .B0(N7375));
XNOR2X1 inst_cellmath__24_0_I2103 (.Y(inst_cellmath__24_0_out0[19]), .A(N2287), .B(N2290));
XNOR2X1 inst_cellmath__24_0_I2104 (.Y(inst_cellmath__24_0_out0[20]), .A(N2349), .B(N2292));
XNOR2X1 inst_cellmath__24_0_I2105 (.Y(inst_cellmath__24_0_out0[21]), .A(N2355), .B(N2294));
XNOR2X1 inst_cellmath__24_0_I2106 (.Y(inst_cellmath__24_0_out0[22]), .A(N2363), .B(N2296));
XNOR2X1 inst_cellmath__24_0_I2107 (.Y(inst_cellmath__24_0_out0[23]), .A(N2373), .B(N2298));
XNOR2X1 inst_cellmath__24_0_I2108 (.Y(inst_cellmath__24_0_out0[24]), .A(N2385), .B(N2300));
XNOR2X1 inst_cellmath__24_0_I2109 (.Y(inst_cellmath__24_0_out0[25]), .A(N2399), .B(N2302));
XNOR2X1 inst_cellmath__24_0_I2110 (.Y(inst_cellmath__24_0_out0[26]), .A(N2415), .B(N2304));
XNOR2X1 inst_cellmath__24_0_I2111 (.Y(inst_cellmath__24_0_out0[27]), .A(N2433), .B(N2306));
XNOR2X1 inst_cellmath__24_0_I2112 (.Y(inst_cellmath__24_0_out0[28]), .A(N2453), .B(N2308));
XNOR2X1 inst_cellmath__24_0_I2113 (.Y(inst_cellmath__24_0_out0[29]), .A(N2475), .B(N2310));
XNOR2X1 inst_cellmath__24_0_I2114 (.Y(inst_cellmath__24_0_out0[30]), .A(N2499), .B(N2312));
XNOR2X1 inst_cellmath__24_0_I2115 (.Y(inst_cellmath__24_0_out0[31]), .A(N2525), .B(N2314));
XNOR2X1 inst_cellmath__24_0_I2116 (.Y(inst_cellmath__24_0_out0[32]), .A(N2553), .B(N2316));
XNOR2X1 inst_cellmath__24_0_I2117 (.Y(inst_cellmath__24_0_out0[33]), .A(N2583), .B(N2318));
XNOR2X1 inst_cellmath__24_0_I2118 (.Y(inst_cellmath__24_0_out0[34]), .A(N2615), .B(N2320));
XNOR2X1 inst_cellmath__24_0_I2119 (.Y(inst_cellmath__24_0_out0[35]), .A(N2649), .B(N2322));
XNOR2X1 inst_cellmath__24_0_I2120 (.Y(inst_cellmath__24_0_out0[36]), .A(N2685), .B(N2324));
XNOR2X1 inst_cellmath__24_0_I2121 (.Y(inst_cellmath__24_0_out0[37]), .A(N2723), .B(N2326));
XNOR2X1 inst_cellmath__24_0_I2122 (.Y(inst_cellmath__24_0_out0[38]), .A(N2763), .B(N2328));
XNOR2X1 inst_cellmath__24_0_I2123 (.Y(inst_cellmath__24_0_out0[39]), .A(N2805), .B(N2330));
XNOR2X1 inst_cellmath__24_0_I2124 (.Y(inst_cellmath__24_0_out0[40]), .A(N2849), .B(N2332));
XNOR2X1 inst_cellmath__24_0_I2125 (.Y(inst_cellmath__24_0_out0[41]), .A(N2895), .B(N2334));
XNOR2X1 inst_cellmath__24_0_I2126 (.Y(inst_cellmath__24_0_out0[42]), .A(N2943), .B(N2336));
XNOR2X1 inst_cellmath__24_0_I2127 (.Y(inst_cellmath__24_0_out0[43]), .A(N2993), .B(N2338));
XNOR2X1 inst_cellmath__24_0_I2128 (.Y(inst_cellmath__24_0_out0[44]), .A(N3045), .B(N2340));
XNOR2X1 inst_cellmath__24_0_I2129 (.Y(inst_cellmath__24_0_out0[45]), .A(N3099), .B(N2342));
XNOR2X1 inst_cellmath__24_0_I2130 (.Y(inst_cellmath__24_0_out0[46]), .A(N3155), .B(N2344));
XOR2XL inst_cellmath__24_0_I3555 (.Y(inst_cellmath__24_0_out0[47]), .A(N3213), .B(N2346));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__25_0_bdw2876250654_bdw (
	inst_cellmath__25_0_out0,
	inst_cellmath__25_0_in0
	); /* architecture "gate_level" */ 
output [47:0] inst_cellmath__25_0_out0;
input [47:0] inst_cellmath__25_0_in0;
wire N199;
BUFX2 inst_cellmath__25_0_I51 (.Y(N199), .A(inst_cellmath__25_0_in0[47]));
AND2XL inst_cellmath__25_0_I0 (.Y(inst_cellmath__25_0_out0[0]), .A(N199), .B(inst_cellmath__25_0_in0[0]));
MX2XL inst_cellmath__25_0_I1 (.Y(inst_cellmath__25_0_out0[1]), .A(inst_cellmath__25_0_in0[0]), .B(inst_cellmath__25_0_in0[1]), .S0(N199));
MX2XL inst_cellmath__25_0_I2 (.Y(inst_cellmath__25_0_out0[2]), .A(inst_cellmath__25_0_in0[1]), .B(inst_cellmath__25_0_in0[2]), .S0(N199));
MX2XL inst_cellmath__25_0_I3 (.Y(inst_cellmath__25_0_out0[3]), .A(inst_cellmath__25_0_in0[2]), .B(inst_cellmath__25_0_in0[3]), .S0(N199));
MX2XL inst_cellmath__25_0_I4 (.Y(inst_cellmath__25_0_out0[4]), .A(inst_cellmath__25_0_in0[3]), .B(inst_cellmath__25_0_in0[4]), .S0(N199));
MX2XL inst_cellmath__25_0_I5 (.Y(inst_cellmath__25_0_out0[5]), .A(inst_cellmath__25_0_in0[4]), .B(inst_cellmath__25_0_in0[5]), .S0(N199));
MX2XL inst_cellmath__25_0_I6 (.Y(inst_cellmath__25_0_out0[6]), .A(inst_cellmath__25_0_in0[5]), .B(inst_cellmath__25_0_in0[6]), .S0(N199));
MX2XL inst_cellmath__25_0_I7 (.Y(inst_cellmath__25_0_out0[7]), .A(inst_cellmath__25_0_in0[6]), .B(inst_cellmath__25_0_in0[7]), .S0(N199));
MX2XL inst_cellmath__25_0_I8 (.Y(inst_cellmath__25_0_out0[8]), .A(inst_cellmath__25_0_in0[7]), .B(inst_cellmath__25_0_in0[8]), .S0(N199));
MX2XL inst_cellmath__25_0_I9 (.Y(inst_cellmath__25_0_out0[9]), .A(inst_cellmath__25_0_in0[8]), .B(inst_cellmath__25_0_in0[9]), .S0(N199));
MX2XL inst_cellmath__25_0_I10 (.Y(inst_cellmath__25_0_out0[10]), .A(inst_cellmath__25_0_in0[9]), .B(inst_cellmath__25_0_in0[10]), .S0(N199));
MX2XL inst_cellmath__25_0_I11 (.Y(inst_cellmath__25_0_out0[11]), .A(inst_cellmath__25_0_in0[10]), .B(inst_cellmath__25_0_in0[11]), .S0(N199));
MX2XL inst_cellmath__25_0_I12 (.Y(inst_cellmath__25_0_out0[12]), .A(inst_cellmath__25_0_in0[11]), .B(inst_cellmath__25_0_in0[12]), .S0(N199));
MX2XL inst_cellmath__25_0_I13 (.Y(inst_cellmath__25_0_out0[13]), .A(inst_cellmath__25_0_in0[12]), .B(inst_cellmath__25_0_in0[13]), .S0(N199));
MX2XL inst_cellmath__25_0_I14 (.Y(inst_cellmath__25_0_out0[14]), .A(inst_cellmath__25_0_in0[13]), .B(inst_cellmath__25_0_in0[14]), .S0(N199));
MX2XL inst_cellmath__25_0_I15 (.Y(inst_cellmath__25_0_out0[15]), .A(inst_cellmath__25_0_in0[14]), .B(inst_cellmath__25_0_in0[15]), .S0(N199));
MX2XL inst_cellmath__25_0_I16 (.Y(inst_cellmath__25_0_out0[16]), .A(inst_cellmath__25_0_in0[15]), .B(inst_cellmath__25_0_in0[16]), .S0(N199));
MX2XL inst_cellmath__25_0_I17 (.Y(inst_cellmath__25_0_out0[17]), .A(inst_cellmath__25_0_in0[16]), .B(inst_cellmath__25_0_in0[17]), .S0(N199));
MX2XL inst_cellmath__25_0_I18 (.Y(inst_cellmath__25_0_out0[18]), .A(inst_cellmath__25_0_in0[17]), .B(inst_cellmath__25_0_in0[18]), .S0(N199));
MX2XL inst_cellmath__25_0_I19 (.Y(inst_cellmath__25_0_out0[19]), .A(inst_cellmath__25_0_in0[18]), .B(inst_cellmath__25_0_in0[19]), .S0(N199));
MX2XL inst_cellmath__25_0_I20 (.Y(inst_cellmath__25_0_out0[20]), .A(inst_cellmath__25_0_in0[19]), .B(inst_cellmath__25_0_in0[20]), .S0(N199));
MX2XL inst_cellmath__25_0_I21 (.Y(inst_cellmath__25_0_out0[21]), .A(inst_cellmath__25_0_in0[20]), .B(inst_cellmath__25_0_in0[21]), .S0(N199));
MX2XL inst_cellmath__25_0_I22 (.Y(inst_cellmath__25_0_out0[22]), .A(inst_cellmath__25_0_in0[21]), .B(inst_cellmath__25_0_in0[22]), .S0(N199));
MX2XL inst_cellmath__25_0_I23 (.Y(inst_cellmath__25_0_out0[23]), .A(inst_cellmath__25_0_in0[22]), .B(inst_cellmath__25_0_in0[23]), .S0(N199));
MX2XL inst_cellmath__25_0_I24 (.Y(inst_cellmath__25_0_out0[24]), .A(inst_cellmath__25_0_in0[23]), .B(inst_cellmath__25_0_in0[24]), .S0(N199));
MX2XL inst_cellmath__25_0_I25 (.Y(inst_cellmath__25_0_out0[25]), .A(inst_cellmath__25_0_in0[24]), .B(inst_cellmath__25_0_in0[25]), .S0(N199));
MX2XL inst_cellmath__25_0_I26 (.Y(inst_cellmath__25_0_out0[26]), .A(inst_cellmath__25_0_in0[25]), .B(inst_cellmath__25_0_in0[26]), .S0(N199));
MX2XL inst_cellmath__25_0_I27 (.Y(inst_cellmath__25_0_out0[27]), .A(inst_cellmath__25_0_in0[26]), .B(inst_cellmath__25_0_in0[27]), .S0(N199));
MX2XL inst_cellmath__25_0_I28 (.Y(inst_cellmath__25_0_out0[28]), .A(inst_cellmath__25_0_in0[27]), .B(inst_cellmath__25_0_in0[28]), .S0(N199));
MX2XL inst_cellmath__25_0_I29 (.Y(inst_cellmath__25_0_out0[29]), .A(inst_cellmath__25_0_in0[28]), .B(inst_cellmath__25_0_in0[29]), .S0(N199));
MX2XL inst_cellmath__25_0_I30 (.Y(inst_cellmath__25_0_out0[30]), .A(inst_cellmath__25_0_in0[29]), .B(inst_cellmath__25_0_in0[30]), .S0(N199));
MX2XL inst_cellmath__25_0_I31 (.Y(inst_cellmath__25_0_out0[31]), .A(inst_cellmath__25_0_in0[30]), .B(inst_cellmath__25_0_in0[31]), .S0(N199));
MX2XL inst_cellmath__25_0_I32 (.Y(inst_cellmath__25_0_out0[32]), .A(inst_cellmath__25_0_in0[31]), .B(inst_cellmath__25_0_in0[32]), .S0(N199));
MX2XL inst_cellmath__25_0_I33 (.Y(inst_cellmath__25_0_out0[33]), .A(inst_cellmath__25_0_in0[32]), .B(inst_cellmath__25_0_in0[33]), .S0(N199));
MX2XL inst_cellmath__25_0_I34 (.Y(inst_cellmath__25_0_out0[34]), .A(inst_cellmath__25_0_in0[33]), .B(inst_cellmath__25_0_in0[34]), .S0(N199));
MX2XL inst_cellmath__25_0_I35 (.Y(inst_cellmath__25_0_out0[35]), .A(inst_cellmath__25_0_in0[34]), .B(inst_cellmath__25_0_in0[35]), .S0(N199));
MX2XL inst_cellmath__25_0_I36 (.Y(inst_cellmath__25_0_out0[36]), .A(inst_cellmath__25_0_in0[35]), .B(inst_cellmath__25_0_in0[36]), .S0(N199));
MX2XL inst_cellmath__25_0_I37 (.Y(inst_cellmath__25_0_out0[37]), .A(inst_cellmath__25_0_in0[36]), .B(inst_cellmath__25_0_in0[37]), .S0(N199));
MX2XL inst_cellmath__25_0_I38 (.Y(inst_cellmath__25_0_out0[38]), .A(inst_cellmath__25_0_in0[37]), .B(inst_cellmath__25_0_in0[38]), .S0(N199));
MX2XL inst_cellmath__25_0_I39 (.Y(inst_cellmath__25_0_out0[39]), .A(inst_cellmath__25_0_in0[38]), .B(inst_cellmath__25_0_in0[39]), .S0(N199));
MX2XL inst_cellmath__25_0_I40 (.Y(inst_cellmath__25_0_out0[40]), .A(inst_cellmath__25_0_in0[39]), .B(inst_cellmath__25_0_in0[40]), .S0(N199));
MX2XL inst_cellmath__25_0_I41 (.Y(inst_cellmath__25_0_out0[41]), .A(inst_cellmath__25_0_in0[40]), .B(inst_cellmath__25_0_in0[41]), .S0(N199));
MX2XL inst_cellmath__25_0_I42 (.Y(inst_cellmath__25_0_out0[42]), .A(inst_cellmath__25_0_in0[41]), .B(inst_cellmath__25_0_in0[42]), .S0(N199));
MX2XL inst_cellmath__25_0_I43 (.Y(inst_cellmath__25_0_out0[43]), .A(inst_cellmath__25_0_in0[42]), .B(inst_cellmath__25_0_in0[43]), .S0(N199));
MX2XL inst_cellmath__25_0_I44 (.Y(inst_cellmath__25_0_out0[44]), .A(inst_cellmath__25_0_in0[43]), .B(inst_cellmath__25_0_in0[44]), .S0(N199));
MX2XL inst_cellmath__25_0_I45 (.Y(inst_cellmath__25_0_out0[45]), .A(inst_cellmath__25_0_in0[44]), .B(inst_cellmath__25_0_in0[45]), .S0(N199));
MX2XL inst_cellmath__25_0_I46 (.Y(inst_cellmath__25_0_out0[46]), .A(inst_cellmath__25_0_in0[45]), .B(inst_cellmath__25_0_in0[46]), .S0(N199));
OR2XL inst_cellmath__25_0_I47 (.Y(inst_cellmath__25_0_out0[47]), .A(N199), .B(inst_cellmath__25_0_in0[46]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__45_0_bdw2876250654_bdw (
	inst_cellmath__45_0_out0,
	inst_cellmath__45_0_in0
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__45_0_out0;
input [47:24] inst_cellmath__45_0_in0;
wire N146,N154,N160,N164,N172,N181,N184 
	,N187,N190,N196,N200,N208,N212,N216,N224 
	,N238,N240,N263,N272,N278,N284,N288,N296 
	,N300,N312,N328,N348,N381,N384,N387,N390 
	,N393,N396,N399,N402,N733,N743,N749,N750 
	,N752,N753,N755,N763;
INVXL inst_cellmath__45_0_I37 (.Y(inst_cellmath__45_0_out0[0]), .A(inst_cellmath__45_0_in0[24]));
NAND2XL inst_cellmath__45_0_I42 (.Y(N146), .A(inst_cellmath__45_0_in0[26]), .B(inst_cellmath__45_0_in0[25]));
NOR2X1 inst_cellmath__45_0_I49 (.Y(N154), .A(N146), .B(inst_cellmath__45_0_out0[0]));
NAND2XL inst_cellmath__45_0_I54 (.Y(N160), .A(inst_cellmath__45_0_in0[28]), .B(inst_cellmath__45_0_in0[27]));
NAND2XL inst_cellmath__45_0_I58 (.Y(N164), .A(inst_cellmath__45_0_in0[30]), .B(inst_cellmath__45_0_in0[29]));
NOR2XL inst_cellmath__45_0_I66 (.Y(N172), .A(N164), .B(N160));
NAND2XL inst_cellmath__45_0_I75 (.Y(N181), .A(inst_cellmath__45_0_in0[27]), .B(N154));
NAND2BXL inst_cellmath__45_0_I565 (.Y(N184), .AN(N160), .B(N154));
NAND3BXL inst_cellmath__45_0_I566 (.Y(N187), .AN(N160), .B(inst_cellmath__45_0_in0[29]), .C(N154));
NAND2X2 inst_cellmath__45_0_I81 (.Y(N190), .A(N172), .B(N154));
NAND2XL inst_cellmath__45_0_I86 (.Y(N196), .A(inst_cellmath__45_0_in0[32]), .B(inst_cellmath__45_0_in0[31]));
NAND2XL inst_cellmath__45_0_I90 (.Y(N200), .A(inst_cellmath__45_0_in0[34]), .B(inst_cellmath__45_0_in0[33]));
NOR2XL inst_cellmath__45_0_I98 (.Y(N208), .A(N200), .B(N196));
NAND2XL inst_cellmath__45_0_I102 (.Y(N212), .A(inst_cellmath__45_0_in0[36]), .B(inst_cellmath__45_0_in0[35]));
NAND2XL inst_cellmath__45_0_I106 (.Y(N216), .A(inst_cellmath__45_0_in0[38]), .B(inst_cellmath__45_0_in0[37]));
NOR2XL inst_cellmath__45_0_I114 (.Y(N224), .A(N216), .B(N212));
NAND3BXL inst_cellmath__45_0_I575 (.Y(N238), .AN(N212), .B(inst_cellmath__45_0_in0[37]), .C(N208));
NAND2X1 inst_cellmath__45_0_I130 (.Y(N240), .A(N224), .B(N208));
NOR3BXL inst_cellmath__45_0_I577 (.Y(N263), .AN(inst_cellmath__45_0_in0[33]), .B(N196), .C(N190));
NOR3BXL inst_cellmath__45_0_I579 (.Y(N272), .AN(N208), .B(N212), .C(N190));
NOR2X2 inst_cellmath__45_0_I161 (.Y(N278), .A(N240), .B(N190));
NAND2XL inst_cellmath__45_0_I166 (.Y(N284), .A(inst_cellmath__45_0_in0[40]), .B(inst_cellmath__45_0_in0[39]));
NAND2XL inst_cellmath__45_0_I170 (.Y(N288), .A(inst_cellmath__45_0_in0[42]), .B(inst_cellmath__45_0_in0[41]));
NOR2XL inst_cellmath__45_0_I178 (.Y(N296), .A(N288), .B(N284));
NAND2XL inst_cellmath__45_0_I182 (.Y(N300), .A(inst_cellmath__45_0_in0[44]), .B(inst_cellmath__45_0_in0[43]));
NAND2XL hyperpropagate_3_1_A_I627 (.Y(N763), .A(inst_cellmath__45_0_in0[46]), .B(inst_cellmath__45_0_in0[45]));
NOR2XL hyperpropagate_3_1_A_I628 (.Y(N312), .A(N300), .B(N763));
NAND2XL inst_cellmath__45_0_I210 (.Y(N328), .A(N312), .B(N296));
INVXL inst_cellmath__45_0_I531 (.Y(N733), .A(inst_cellmath__45_0_in0[47]));
NOR2XL inst_cellmath__45_0_I230 (.Y(N348), .A(N733), .B(N328));
NAND2BXL inst_cellmath__45_0_I593 (.Y(N743), .AN(inst_cellmath__45_0_out0[0]), .B(inst_cellmath__45_0_in0[25]));
NAND2BXL inst_cellmath__45_0_I594 (.Y(N749), .AN(N190), .B(inst_cellmath__45_0_in0[31]));
OR2XL inst_cellmath__45_0_I595 (.Y(N750), .A(N196), .B(N190));
NAND2BXL inst_cellmath__45_0_I596 (.Y(N752), .AN(N190), .B(N208));
NAND3BXL inst_cellmath__45_0_I616 (.Y(N753), .AN(N190), .B(inst_cellmath__45_0_in0[35]), .C(N208));
OR2XL inst_cellmath__45_0_I598 (.Y(N755), .A(N238), .B(N190));
NAND2XL inst_cellmath__45_0_I263 (.Y(N381), .A(inst_cellmath__45_0_in0[39]), .B(N278));
NAND2BXL inst_cellmath__45_0_I599 (.Y(N384), .AN(N284), .B(N278));
NAND3BXL inst_cellmath__45_0_I600 (.Y(N387), .AN(N284), .B(inst_cellmath__45_0_in0[41]), .C(N278));
NAND2XL inst_cellmath__45_0_I269 (.Y(N390), .A(N296), .B(N278));
NAND3XL inst_cellmath__45_0_I601 (.Y(N393), .A(inst_cellmath__45_0_in0[43]), .B(N296), .C(N278));
NAND3BXL inst_cellmath__45_0_I602 (.Y(N396), .AN(N300), .B(N296), .C(N278));
NAND4BXL inst_cellmath__45_0_I603 (.Y(N399), .AN(N300), .B(inst_cellmath__45_0_in0[45]), .C(N278), .D(N296));
NAND2BXL inst_cellmath__45_0_I604 (.Y(N402), .AN(N328), .B(N278));
AND2XL inst_cellmath__45_0_I279 (.Y(inst_cellmath__45_0_out0[24]), .A(N348), .B(N278));
XNOR2X1 inst_cellmath__45_0_I380 (.Y(inst_cellmath__45_0_out0[1]), .A(inst_cellmath__45_0_out0[0]), .B(inst_cellmath__45_0_in0[25]));
XNOR2X1 inst_cellmath__45_0_I381 (.Y(inst_cellmath__45_0_out0[2]), .A(N743), .B(inst_cellmath__45_0_in0[26]));
XOR2XL inst_cellmath__45_0_I606 (.Y(inst_cellmath__45_0_out0[3]), .A(N154), .B(inst_cellmath__45_0_in0[27]));
XNOR2X1 inst_cellmath__45_0_I383 (.Y(inst_cellmath__45_0_out0[4]), .A(N181), .B(inst_cellmath__45_0_in0[28]));
XNOR2X1 inst_cellmath__45_0_I384 (.Y(inst_cellmath__45_0_out0[5]), .A(N184), .B(inst_cellmath__45_0_in0[29]));
XNOR2X1 inst_cellmath__45_0_I385 (.Y(inst_cellmath__45_0_out0[6]), .A(N187), .B(inst_cellmath__45_0_in0[30]));
XNOR2X1 inst_cellmath__45_0_I386 (.Y(inst_cellmath__45_0_out0[7]), .A(N190), .B(inst_cellmath__45_0_in0[31]));
XNOR2X1 inst_cellmath__45_0_I387 (.Y(inst_cellmath__45_0_out0[8]), .A(N749), .B(inst_cellmath__45_0_in0[32]));
XNOR2X1 inst_cellmath__45_0_I388 (.Y(inst_cellmath__45_0_out0[9]), .A(N750), .B(inst_cellmath__45_0_in0[33]));
XOR2XL inst_cellmath__45_0_I607 (.Y(inst_cellmath__45_0_out0[10]), .A(N263), .B(inst_cellmath__45_0_in0[34]));
XNOR2X1 inst_cellmath__45_0_I390 (.Y(inst_cellmath__45_0_out0[11]), .A(N752), .B(inst_cellmath__45_0_in0[35]));
XNOR2X1 inst_cellmath__45_0_I391 (.Y(inst_cellmath__45_0_out0[12]), .A(N753), .B(inst_cellmath__45_0_in0[36]));
XOR2XL inst_cellmath__45_0_I608 (.Y(inst_cellmath__45_0_out0[13]), .A(N272), .B(inst_cellmath__45_0_in0[37]));
XNOR2X1 inst_cellmath__45_0_I393 (.Y(inst_cellmath__45_0_out0[14]), .A(N755), .B(inst_cellmath__45_0_in0[38]));
XOR2XL inst_cellmath__45_0_I609 (.Y(inst_cellmath__45_0_out0[15]), .A(N278), .B(inst_cellmath__45_0_in0[39]));
XNOR2X1 inst_cellmath__45_0_I395 (.Y(inst_cellmath__45_0_out0[16]), .A(N381), .B(inst_cellmath__45_0_in0[40]));
XNOR2X1 inst_cellmath__45_0_I396 (.Y(inst_cellmath__45_0_out0[17]), .A(N384), .B(inst_cellmath__45_0_in0[41]));
XNOR2X1 inst_cellmath__45_0_I397 (.Y(inst_cellmath__45_0_out0[18]), .A(N387), .B(inst_cellmath__45_0_in0[42]));
XNOR2X1 inst_cellmath__45_0_I398 (.Y(inst_cellmath__45_0_out0[19]), .A(N390), .B(inst_cellmath__45_0_in0[43]));
XNOR2X1 inst_cellmath__45_0_I399 (.Y(inst_cellmath__45_0_out0[20]), .A(N393), .B(inst_cellmath__45_0_in0[44]));
XNOR2X1 inst_cellmath__45_0_I400 (.Y(inst_cellmath__45_0_out0[21]), .A(N396), .B(inst_cellmath__45_0_in0[45]));
XNOR2X1 inst_cellmath__45_0_I401 (.Y(inst_cellmath__45_0_out0[22]), .A(N399), .B(inst_cellmath__45_0_in0[46]));
XOR2XL inst_cellmath__45_0_I610 (.Y(inst_cellmath__45_0_out0[23]), .A(N733), .B(N402));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__5_1_bdw2876250654_bdw (
	inst_cellmath__5_1_out0,
	inst_cellmath__5_1_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__5_1_out0;
input [2:0] inst_cellmath__5_1_in0;
NOR3BXL inst_cellmath__5_1_I17 (.Y(inst_cellmath__5_1_out0), .AN(inst_cellmath__5_1_in0[0]), .B(inst_cellmath__5_1_in0[2]), .C(inst_cellmath__5_1_in0[1]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__31__bdw2876250654_bdw (
	inst_cellmath__44__31__out0,
	inst_cellmath__44__31__in0,
	inst_cellmath__44__31__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__31__out0;
input  inst_cellmath__44__31__in0,
	inst_cellmath__44__31__in1;
wire N13;
INVXL inst_cellmath__44__31__I3 (.Y(N13), .A(inst_cellmath__44__31__in1));
AND2XL inst_cellmath__44__31__I1 (.Y(inst_cellmath__44__31__out0[0]), .A(inst_cellmath__44__31__in0), .B(N13));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__6_0_bdw2876250654_bdw (
	inst_cellmath__6_0_out0,
	inst_cellmath__6_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__6_0_out0;
input [2:0] inst_cellmath__6_0_in0;
NOR3BXL inst_cellmath__6_0_I23 (.Y(inst_cellmath__6_0_out0), .AN(inst_cellmath__6_0_in0[1]), .B(inst_cellmath__6_0_in0[2]), .C(inst_cellmath__6_0_in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__30__bdw2876250654_bdw (
	inst_cellmath__44__30__out0,
	inst_cellmath__44__30__in0,
	inst_cellmath__44__30__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__30__out0;
input  inst_cellmath__44__30__in0,
	inst_cellmath__44__30__in1;
AND2XL inst_cellmath__44__30__I0 (.Y(inst_cellmath__44__30__out0[0]), .A(inst_cellmath__44__30__in0), .B(inst_cellmath__44__30__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__8_0_bdw2876250654_bdw (
	inst_cellmath__8_0_out0,
	inst_cellmath__8_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__8_0_out0;
input [2:0] inst_cellmath__8_0_in0;
NOR3BXL inst_cellmath__8_0_I34 (.Y(inst_cellmath__8_0_out0), .AN(inst_cellmath__8_0_in0[2]), .B(inst_cellmath__8_0_in0[1]), .C(inst_cellmath__8_0_in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__4_0_bdw2876250654_bdw (
	inst_cellmath__4_0_out0,
	inst_cellmath__4_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__4_0_out0;
input [2:0] inst_cellmath__4_0_in0;
NOR3XL inst_cellmath__4_0_I39 (.Y(inst_cellmath__4_0_out0), .A(inst_cellmath__4_0_in0[1]), .B(inst_cellmath__4_0_in0[2]), .C(inst_cellmath__4_0_in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__34_0_bdw2876250654_bdw (
	inst_cellmath__34_0_out0,
	inst_cellmath__34_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__34_0_out0;
input [22:0] inst_cellmath__34_0_in0;
wire N29,N30,N31,N32,N33,N34,N35 
	,N36,N37,N38,N39,N40,N42,N43,N45 
	,N48,N49,N70;
NOR2XL inst_cellmath__34_0_I3 (.Y(N29), .A(inst_cellmath__34_0_in0[19]), .B(inst_cellmath__34_0_in0[17]));
NOR2XL inst_cellmath__34_0_I4 (.Y(N30), .A(inst_cellmath__34_0_in0[15]), .B(inst_cellmath__34_0_in0[13]));
NOR2XL inst_cellmath__34_0_I5 (.Y(N31), .A(inst_cellmath__34_0_in0[11]), .B(inst_cellmath__34_0_in0[9]));
NOR2XL inst_cellmath__34_0_I6 (.Y(N32), .A(inst_cellmath__34_0_in0[7]), .B(inst_cellmath__34_0_in0[5]));
NOR2XL inst_cellmath__34_0_I7 (.Y(N33), .A(inst_cellmath__34_0_in0[3]), .B(inst_cellmath__34_0_in0[22]));
NOR2XL inst_cellmath__34_0_I8 (.Y(N34), .A(inst_cellmath__34_0_in0[20]), .B(inst_cellmath__34_0_in0[18]));
NOR2XL inst_cellmath__34_0_I9 (.Y(N35), .A(inst_cellmath__34_0_in0[16]), .B(inst_cellmath__34_0_in0[14]));
NOR2XL inst_cellmath__34_0_I10 (.Y(N36), .A(inst_cellmath__34_0_in0[12]), .B(inst_cellmath__34_0_in0[10]));
NOR2XL inst_cellmath__34_0_I11 (.Y(N37), .A(inst_cellmath__34_0_in0[8]), .B(inst_cellmath__34_0_in0[6]));
NOR2XL inst_cellmath__34_0_I12 (.Y(N38), .A(inst_cellmath__34_0_in0[4]), .B(inst_cellmath__34_0_in0[2]));
NAND2XL inst_cellmath__34_0_I13 (.Y(N39), .A(N29), .B(N30));
NAND2XL inst_cellmath__34_0_I14 (.Y(N40), .A(N31), .B(N32));
NAND2XL inst_cellmath__34_0_I16 (.Y(N42), .A(N35), .B(N36));
NAND2XL inst_cellmath__34_0_I17 (.Y(N43), .A(N37), .B(N38));
NOR4X1 inst_cellmath__34_0_I27 (.Y(N45), .A(inst_cellmath__34_0_in0[0]), .B(inst_cellmath__34_0_in0[1]), .C(inst_cellmath__34_0_in0[21]), .D(N39));
NOR2XL inst_cellmath__34_0_I21 (.Y(N49), .A(N42), .B(N43));
NAND3XL hyperpropagate_4_1_A_I30 (.Y(N70), .A(N33), .B(N34), .C(N45));
NOR2XL hyperpropagate_4_1_A_I31 (.Y(N48), .A(N40), .B(N70));
NAND2X1 inst_cellmath__34_0_I24 (.Y(inst_cellmath__34_0_out0), .A(N49), .B(N48));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__29__bdw2876250654_bdw (
	inst_cellmath__44__29__out0,
	inst_cellmath__44__29__in0,
	inst_cellmath__44__29__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__29__out0;
input  inst_cellmath__44__29__in0;
input [24:24] inst_cellmath__44__29__in1;
OR2XL inst_cellmath__44__29__I0 (.Y(inst_cellmath__44__29__out0[0]), .A(inst_cellmath__44__29__in1[24]), .B(inst_cellmath__44__29__in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__28__bdw2876250654_bdw (
	inst_cellmath__44__28__out0,
	inst_cellmath__44__28__in0,
	inst_cellmath__44__28__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__28__out0;
input [0:0] inst_cellmath__44__28__in0;
input  inst_cellmath__44__28__in1;
AND2XL inst_cellmath__44__28__I0 (.Y(inst_cellmath__44__28__out0[0]), .A(inst_cellmath__44__28__in1), .B(inst_cellmath__44__28__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__27__bdw2876250654_bdw (
	inst_cellmath__44__27__out0,
	inst_cellmath__44__27__in0,
	inst_cellmath__44__27__in1,
	inst_cellmath__44__27__in2,
	inst_cellmath__44__27__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__27__out0;
input  inst_cellmath__44__27__in0;
input [0:0] inst_cellmath__44__27__in1,
	inst_cellmath__44__27__in2,
	inst_cellmath__44__27__in3;
OR4X1 inst_cellmath__44__27__I7 (.Y(inst_cellmath__44__27__out0[0]), .A(inst_cellmath__44__27__in0), .B(inst_cellmath__44__27__in2[0]), .C(inst_cellmath__44__27__in1[0]), .D(inst_cellmath__44__27__in3[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__26__bdw2876250654_bdw (
	inst_cellmath__44__26__out0,
	inst_cellmath__44__26__in0,
	inst_cellmath__44__26__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__26__out0;
input [0:0] inst_cellmath__44__26__in0;
input [23:23] inst_cellmath__44__26__in1;
AND2XL inst_cellmath__44__26__I0 (.Y(inst_cellmath__44__26__out0[0]), .A(inst_cellmath__44__26__in1[23]), .B(inst_cellmath__44__26__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__33__bdw2876250654_bdw (
	inst_cellmath__44__33__out0,
	inst_cellmath__44__33__in0,
	inst_cellmath__44__33__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__33__out0;
input [0:0] inst_cellmath__44__33__in0,
	inst_cellmath__44__33__in1;
OR2XL inst_cellmath__44__33__I0 (.Y(inst_cellmath__44__33__out0[0]), .A(inst_cellmath__44__33__in1[0]), .B(inst_cellmath__44__33__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__32__bdw2876250654_bdw (
	inst_cellmath__44__32__out0,
	inst_cellmath__44__32__in0,
	inst_cellmath__44__32__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__32__out0;
input [0:0] inst_cellmath__44__32__in0;
input  inst_cellmath__44__32__in1;
AND2XL inst_cellmath__44__32__I0 (.Y(inst_cellmath__44__32__out0[0]), .A(inst_cellmath__44__32__in0[0]), .B(inst_cellmath__44__32__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44_0_bdw2876250654_bdw (
	inst_cellmath__44_0_out0,
	inst_cellmath__44_0_in0,
	inst_cellmath__44_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__44_0_out0;
input [0:0] inst_cellmath__44_0_in0,
	inst_cellmath__44_0_in1;
OR2XL inst_cellmath__44_0_I0 (.Y(inst_cellmath__44_0_out0), .A(inst_cellmath__44_0_in0[0]), .B(inst_cellmath__44_0_in1[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__46_0_bdw2876250654_bdw (
	inst_cellmath__46_0_out0,
	inst_cellmath__46_0_in0,
	inst_cellmath__46_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__46_0_out0;
input [24:24] inst_cellmath__46_0_in0;
input  inst_cellmath__46_0_in1;
AND2XL inst_cellmath__46_0_I0 (.Y(inst_cellmath__46_0_out0), .A(inst_cellmath__46_0_in0[24]), .B(inst_cellmath__46_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__38_0_bdw2876250654_bdw (
	inst_cellmath__38_0_out0,
	inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__38_0_out0;
input  inst_cellmath__38_0_in0;
input [47:47] inst_cellmath__38_0_in1;
OR2XL inst_cellmath__38_0_I0 (.Y(inst_cellmath__38_0_out0), .A(inst_cellmath__38_0_in1[47]), .B(inst_cellmath__38_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__30_0_bdw2876250654_bdw (
	inst_cellmath__30_0_out0,
	inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__30_0_out0;
input [7:0] inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1;
wire N106,N111,N115,N117,N119,N121,N123 
	,N125,N127;
INVXL inst_cellmath__30_0_I40 (.Y(N106), .A(inst_cellmath__30_0_in1[7]));
XNOR2X1 hap1_A_I51 (.Y(inst_cellmath__30_0_out0[0]), .A(inst_cellmath__30_0_in0[0]), .B(inst_cellmath__30_0_in1[0]));
OR2XL hap1_A_I52 (.Y(N111), .A(inst_cellmath__30_0_in0[0]), .B(inst_cellmath__30_0_in1[0]));
ADDFX1 inst_cellmath__30_0_I42 (.CO(N115), .S(inst_cellmath__30_0_out0[1]), .A(inst_cellmath__30_0_in0[1]), .B(inst_cellmath__30_0_in1[1]), .CI(N111));
ADDFX1 inst_cellmath__30_0_I43 (.CO(N117), .S(inst_cellmath__30_0_out0[2]), .A(inst_cellmath__30_0_in0[2]), .B(inst_cellmath__30_0_in1[2]), .CI(N115));
ADDFX1 inst_cellmath__30_0_I44 (.CO(N119), .S(inst_cellmath__30_0_out0[3]), .A(inst_cellmath__30_0_in0[3]), .B(inst_cellmath__30_0_in1[3]), .CI(N117));
ADDFX1 inst_cellmath__30_0_I45 (.CO(N121), .S(inst_cellmath__30_0_out0[4]), .A(inst_cellmath__30_0_in0[4]), .B(inst_cellmath__30_0_in1[4]), .CI(N119));
ADDFX1 inst_cellmath__30_0_I46 (.CO(N123), .S(inst_cellmath__30_0_out0[5]), .A(inst_cellmath__30_0_in0[5]), .B(inst_cellmath__30_0_in1[5]), .CI(N121));
ADDFX1 inst_cellmath__30_0_I47 (.CO(N125), .S(inst_cellmath__30_0_out0[6]), .A(inst_cellmath__30_0_in0[6]), .B(inst_cellmath__30_0_in1[6]), .CI(N123));
ADDFX1 inst_cellmath__30_0_I48 (.CO(N127), .S(inst_cellmath__30_0_out0[7]), .A(N106), .B(inst_cellmath__30_0_in0[7]), .CI(N125));
XNOR2X1 hap1_A_I53 (.Y(inst_cellmath__30_0_out0[8]), .A(inst_cellmath__30_0_in1[7]), .B(N127));
NOR2XL hap1_A_I54 (.Y(inst_cellmath__30_0_out0[9]), .A(inst_cellmath__30_0_in1[7]), .B(N127));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__31_0_bdw2876250654_bdw (
	inst_cellmath__31_0_out0,
	inst_cellmath__31_0_in0
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__31_0_out0;
input [9:0] inst_cellmath__31_0_in0;
wire N77,N116,N119,N128,N131,N134,N137 
	,N140;
INVXL inst_cellmath__31_0_I99 (.Y(inst_cellmath__31_0_out0[0]), .A(inst_cellmath__31_0_in0[0]));
NOR2BX1 inst_cellmath__31_0_I102 (.Y(N77), .AN(inst_cellmath__31_0_in0[1]), .B(inst_cellmath__31_0_out0[0]));
AND2XL inst_cellmath__31_0_I38 (.Y(N116), .A(inst_cellmath__31_0_in0[2]), .B(N77));
XNOR2X1 inst_cellmath__31_0_I55 (.Y(inst_cellmath__31_0_out0[1]), .A(inst_cellmath__31_0_out0[0]), .B(inst_cellmath__31_0_in0[1]));
XOR2XL inst_cellmath__31_0_I103 (.Y(inst_cellmath__31_0_out0[2]), .A(N77), .B(inst_cellmath__31_0_in0[2]));
AND2XL inst_cellmath__31_0_I60 (.Y(N119), .A(inst_cellmath__31_0_in0[3]), .B(N116));
AND3XL inst_cellmath__31_0_I104 (.Y(N128), .A(inst_cellmath__31_0_in0[4]), .B(inst_cellmath__31_0_in0[5]), .C(N119));
AND3XL inst_cellmath__31_0_I105 (.Y(N131), .A(inst_cellmath__31_0_in0[6]), .B(inst_cellmath__31_0_in0[7]), .C(N128));
NAND2XL inst_cellmath__31_0_I72 (.Y(N134), .A(inst_cellmath__31_0_in0[4]), .B(N119));
NAND2XL inst_cellmath__31_0_I74 (.Y(N137), .A(inst_cellmath__31_0_in0[6]), .B(N128));
NAND2XL inst_cellmath__31_0_I76 (.Y(N140), .A(inst_cellmath__31_0_in0[8]), .B(N131));
XOR2XL inst_cellmath__31_0_I84 (.Y(inst_cellmath__31_0_out0[3]), .A(N116), .B(inst_cellmath__31_0_in0[3]));
XOR2XL inst_cellmath__31_0_I85 (.Y(inst_cellmath__31_0_out0[4]), .A(N119), .B(inst_cellmath__31_0_in0[4]));
XNOR2X1 inst_cellmath__31_0_I86 (.Y(inst_cellmath__31_0_out0[5]), .A(N134), .B(inst_cellmath__31_0_in0[5]));
XOR2XL inst_cellmath__31_0_I87 (.Y(inst_cellmath__31_0_out0[6]), .A(N128), .B(inst_cellmath__31_0_in0[6]));
XNOR2X1 inst_cellmath__31_0_I88 (.Y(inst_cellmath__31_0_out0[7]), .A(N137), .B(inst_cellmath__31_0_in0[7]));
XOR2XL inst_cellmath__31_0_I89 (.Y(inst_cellmath__31_0_out0[8]), .A(N131), .B(inst_cellmath__31_0_in0[8]));
XNOR2X1 inst_cellmath__31_0_I90 (.Y(inst_cellmath__31_0_out0[9]), .A(N140), .B(inst_cellmath__31_0_in0[9]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__48_0_bdw2876250654_bdw (
	inst_cellmath__48_0_out0,
	inst_cellmath__48_0_in0,
	inst_cellmath__48_0_in1,
	inst_cellmath__48_0_in2
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__48_0_out0;
input  inst_cellmath__48_0_in0;
input [9:0] inst_cellmath__48_0_in1,
	inst_cellmath__48_0_in2;
MX2XL inst_cellmath__48_0_I20 (.Y(inst_cellmath__48_0_out0[0]), .A(inst_cellmath__48_0_in2[0]), .B(inst_cellmath__48_0_in1[0]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I21 (.Y(inst_cellmath__48_0_out0[1]), .A(inst_cellmath__48_0_in2[1]), .B(inst_cellmath__48_0_in1[1]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I22 (.Y(inst_cellmath__48_0_out0[2]), .A(inst_cellmath__48_0_in2[2]), .B(inst_cellmath__48_0_in1[2]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I23 (.Y(inst_cellmath__48_0_out0[3]), .A(inst_cellmath__48_0_in2[3]), .B(inst_cellmath__48_0_in1[3]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I24 (.Y(inst_cellmath__48_0_out0[4]), .A(inst_cellmath__48_0_in2[4]), .B(inst_cellmath__48_0_in1[4]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I25 (.Y(inst_cellmath__48_0_out0[5]), .A(inst_cellmath__48_0_in2[5]), .B(inst_cellmath__48_0_in1[5]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I26 (.Y(inst_cellmath__48_0_out0[6]), .A(inst_cellmath__48_0_in2[6]), .B(inst_cellmath__48_0_in1[6]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I27 (.Y(inst_cellmath__48_0_out0[7]), .A(inst_cellmath__48_0_in2[7]), .B(inst_cellmath__48_0_in1[7]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I28 (.Y(inst_cellmath__48_0_out0[8]), .A(inst_cellmath__48_0_in2[8]), .B(inst_cellmath__48_0_in1[8]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I29 (.Y(inst_cellmath__48_0_out0[9]), .A(inst_cellmath__48_0_in2[9]), .B(inst_cellmath__48_0_in1[9]), .S0(inst_cellmath__48_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51__49__bdw2876250654_bdw (
	inst_cellmath__51__49__out0,
	inst_cellmath__51__49__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__51__49__out0;
input [7:0] inst_cellmath__51__49__in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__51__49__I0 (.Y(N11), .A(inst_cellmath__51__49__in0[1]), .B(inst_cellmath__51__49__in0[6]));
NAND2XL inst_cellmath__51__49__I1 (.Y(N12), .A(inst_cellmath__51__49__in0[0]), .B(inst_cellmath__51__49__in0[5]));
NAND2XL inst_cellmath__51__49__I2 (.Y(N13), .A(inst_cellmath__51__49__in0[4]), .B(inst_cellmath__51__49__in0[2]));
NAND2XL inst_cellmath__51__49__I3 (.Y(N14), .A(inst_cellmath__51__49__in0[7]), .B(inst_cellmath__51__49__in0[3]));
NOR2XL inst_cellmath__51__49__I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__51__49__I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__51__49__I6 (.Y(inst_cellmath__51__49__out0[0]), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51__48__bdw2876250654_bdw (
	inst_cellmath__51__48__out0,
	inst_cellmath__51__48__in0,
	inst_cellmath__51__48__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__51__48__out0;
input [0:0] inst_cellmath__51__48__in0;
input [8:8] inst_cellmath__51__48__in1;
OR2XL inst_cellmath__51__48__I0 (.Y(inst_cellmath__51__48__out0[0]), .A(inst_cellmath__51__48__in1[8]), .B(inst_cellmath__51__48__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51_0_bdw2876250654_bdw (
	inst_cellmath__51_0_out0,
	inst_cellmath__51_0_in0,
	inst_cellmath__51_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__51_0_out0;
input [0:0] inst_cellmath__51_0_in0;
input [9:9] inst_cellmath__51_0_in1;
NOR2BX1 inst_cellmath__51_0_I3 (.Y(inst_cellmath__51_0_out0), .AN(inst_cellmath__51_0_in0[0]), .B(inst_cellmath__51_0_in1[9]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__28_0_bdw2876250654_bdw (
	inst_cellmath__28_0_out0,
	inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__28_0_out0;
input  inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1;
OR2XL inst_cellmath__28_0_I0 (.Y(inst_cellmath__28_0_out0), .A(inst_cellmath__28_0_in0), .B(inst_cellmath__28_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__27_0_bdw2876250654_bdw (
	inst_cellmath__27_0_out0,
	inst_cellmath__27_0_in0,
	inst_cellmath__27_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__27_0_out0;
input  inst_cellmath__27_0_in0,
	inst_cellmath__27_0_in1;
OR2XL inst_cellmath__27_0_I0 (.Y(inst_cellmath__27_0_out0), .A(inst_cellmath__27_0_in0), .B(inst_cellmath__27_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__50__50__bdw2876250654_bdw (
	inst_cellmath__50__50__out0,
	inst_cellmath__50__50__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__50__50__out0;
input [9:0] inst_cellmath__50__50__in0;
wire N13,N14,N18,N21,N22;
NOR2XL inst_cellmath__50__50__I0 (.Y(N13), .A(inst_cellmath__50__50__in0[8]), .B(inst_cellmath__50__50__in0[1]));
NOR2XL inst_cellmath__50__50__I1 (.Y(N14), .A(inst_cellmath__50__50__in0[6]), .B(inst_cellmath__50__50__in0[9]));
NAND2XL inst_cellmath__50__50__I5 (.Y(N18), .A(N13), .B(N14));
NOR4X1 inst_cellmath__50__50__I13 (.Y(N22), .A(inst_cellmath__50__50__in0[0]), .B(inst_cellmath__50__50__in0[2]), .C(inst_cellmath__50__50__in0[4]), .D(inst_cellmath__50__50__in0[5]));
NOR3XL inst_cellmath__50__50__I12 (.Y(N21), .A(inst_cellmath__50__50__in0[7]), .B(inst_cellmath__50__50__in0[3]), .C(N18));
NAND2XL inst_cellmath__50__50__I10 (.Y(inst_cellmath__50__50__out0[0]), .A(N22), .B(N21));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__49_1_bdw2876250654_bdw (
	inst_cellmath__49_1_out0,
	inst_cellmath__49_1_in0,
	inst_cellmath__49_1_in1,
	inst_cellmath__49_1_in2,
	inst_cellmath__49_1_in3,
	inst_cellmath__49_1_in4,
	inst_cellmath__49_1_in5
	); /* architecture "gate_level" */ 
output  inst_cellmath__49_1_out0;
input  inst_cellmath__49_1_in0;
input [0:0] inst_cellmath__49_1_in1;
input [9:9] inst_cellmath__49_1_in2;
input  inst_cellmath__49_1_in3,
	inst_cellmath__49_1_in4,
	inst_cellmath__49_1_in5;
wire N13,N14;
NOR4XL inst_cellmath__49_1_I9 (.Y(N13), .A(inst_cellmath__49_1_in3), .B(inst_cellmath__49_1_in4), .C(inst_cellmath__49_1_in5), .D(inst_cellmath__49_1_in2[9]));
NAND2XL inst_cellmath__49_1_I5 (.Y(N14), .A(N13), .B(inst_cellmath__49_1_in1[0]));
OR2XL inst_cellmath__49_1_I6 (.Y(inst_cellmath__49_1_out0), .A(N14), .B(inst_cellmath__49_1_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__37__43__bdw2876250654_bdw (
	inst_cellmath__37__43__out0,
	inst_cellmath__37__43__in0,
	inst_cellmath__37__43__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__37__43__out0;
input  inst_cellmath__37__43__in0,
	inst_cellmath__37__43__in1;
OR2XL inst_cellmath__37__43__I0 (.Y(inst_cellmath__37__43__out0[0]), .A(inst_cellmath__37__43__in0), .B(inst_cellmath__37__43__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__32__11__bdw2876250654_bdw (
	inst_cellmath__32__11__out0,
	inst_cellmath__32__11__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__32__11__out0;
input [8:7] inst_cellmath__32__11__in0;
OR2XL inst_cellmath__32__11__I0 (.Y(inst_cellmath__32__11__out0[0]), .A(inst_cellmath__32__11__in0[8]), .B(inst_cellmath__32__11__in0[7]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__32__10__bdw2876250654_bdw (
	inst_cellmath__32__10__out0,
	inst_cellmath__32__10__in0,
	inst_cellmath__32__10__in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__32__10__out0;
input [0:0] inst_cellmath__32__10__in0;
input [9:9] inst_cellmath__32__10__in1;
NAND2BXL inst_cellmath__32__10__I2 (.Y(inst_cellmath__32__10__out0), .AN(inst_cellmath__32__10__in1[9]), .B(inst_cellmath__32__10__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__37__42__bdw2876250654_bdw (
	inst_cellmath__37__42__out0,
	inst_cellmath__37__42__in0,
	inst_cellmath__37__42__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__37__42__out0;
input  inst_cellmath__37__42__in0,
	inst_cellmath__37__42__in1;
OR2XL inst_cellmath__37__42__I0 (.Y(inst_cellmath__37__42__out0[0]), .A(inst_cellmath__37__42__in1), .B(inst_cellmath__37__42__in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__7_0_bdw2876250654_bdw (
	inst_cellmath__7_0_out0,
	inst_cellmath__7_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__7_0_out0;
input [2:0] inst_cellmath__7_0_in0;
wire N42;
NAND2XL inst_cellmath__7_0_I24 (.Y(N42), .A(inst_cellmath__7_0_in0[0]), .B(inst_cellmath__7_0_in0[1]));
NOR2XL inst_cellmath__7_0_I25 (.Y(inst_cellmath__7_0_out0), .A(inst_cellmath__7_0_in0[2]), .B(N42));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__42_0_bdw2876250654_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1,
	inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__42_0_out0;
input  inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1,
	inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3;
wire N12,N21;
INVXL inst_cellmath__42_0_I6 (.Y(N21), .A(inst_cellmath__42_0_in3));
MXI2XL inst_cellmath__42_0_I3 (.Y(N12), .A(inst_cellmath__42_0_in0), .B(N21), .S0(inst_cellmath__42_0_in1));
MX2XL inst_cellmath__42_0_I4 (.Y(inst_cellmath__42_0_out0), .A(N12), .B(N21), .S0(inst_cellmath__42_0_in2));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__52_0_bdw2876250654_bdw (
	inst_cellmath__52_0_out0,
	inst_cellmath__52_0_in0,
	inst_cellmath__52_0_in1,
	inst_cellmath__52_0_in2,
	inst_cellmath__52_0_in3,
	inst_cellmath__52_0_in4
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__52_0_out0;
input  inst_cellmath__52_0_in0;
input [7:0] inst_cellmath__52_0_in1;
input  inst_cellmath__52_0_in2;
input [0:0] inst_cellmath__52_0_in3,
	inst_cellmath__52_0_in4;
wire N50,N134,N136,N137,N138,N141;
INVXL inst_cellmath__52_0_I54 (.Y(N137), .A(inst_cellmath__52_0_in4[0]));
AOI21XL inst_cellmath__52_0_I56 (.Y(N50), .A0(inst_cellmath__52_0_in2), .A1(N137), .B0(inst_cellmath__52_0_in3[0]));
OR2XL inst_cellmath__52_0_I57 (.Y(N134), .A(N137), .B(inst_cellmath__52_0_in3[0]));
INVXL inst_cellmath__52_0_I55 (.Y(N138), .A(inst_cellmath__52_0_in1[0]));
INVXL buf1_A_I59 (.Y(N141), .A(inst_cellmath__52_0_in0));
INVXL buf1_A_I60 (.Y(N136), .A(N141));
MXI2XL inst_cellmath__52_0_I32 (.Y(inst_cellmath__52_0_out0[0]), .A(N138), .B(N50), .S0(N136));
MX2XL inst_cellmath__52_0_I33 (.Y(inst_cellmath__52_0_out0[1]), .A(inst_cellmath__52_0_in1[1]), .B(N134), .S0(N136));
MX2XL inst_cellmath__52_0_I34 (.Y(inst_cellmath__52_0_out0[2]), .A(inst_cellmath__52_0_in1[2]), .B(N134), .S0(N136));
MX2XL inst_cellmath__52_0_I35 (.Y(inst_cellmath__52_0_out0[3]), .A(inst_cellmath__52_0_in1[3]), .B(N134), .S0(N136));
MX2XL inst_cellmath__52_0_I36 (.Y(inst_cellmath__52_0_out0[4]), .A(inst_cellmath__52_0_in1[4]), .B(N134), .S0(N136));
MX2XL inst_cellmath__52_0_I37 (.Y(inst_cellmath__52_0_out0[5]), .A(inst_cellmath__52_0_in1[5]), .B(N134), .S0(N136));
MX2XL inst_cellmath__52_0_I38 (.Y(inst_cellmath__52_0_out0[6]), .A(inst_cellmath__52_0_in1[6]), .B(N134), .S0(N136));
MX2XL inst_cellmath__52_0_I39 (.Y(inst_cellmath__52_0_out0[7]), .A(inst_cellmath__52_0_in1[7]), .B(N134), .S0(N136));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__47_0_bdw2876250654_bdw (
	inst_cellmath__47_0_out0,
	inst_cellmath__47_0_in0,
	inst_cellmath__47_0_in1,
	inst_cellmath__47_0_in2,
	inst_cellmath__47_0_in3,
	inst_cellmath__47_0_in4
	); /* architecture "gate_level" */ 
output  inst_cellmath__47_0_out0;
input  inst_cellmath__47_0_in0,
	inst_cellmath__47_0_in1,
	inst_cellmath__47_0_in2,
	inst_cellmath__47_0_in3,
	inst_cellmath__47_0_in4;
wire N12;
OR4X1 inst_cellmath__47_0_I7 (.Y(N12), .A(inst_cellmath__47_0_in2), .B(inst_cellmath__47_0_in3), .C(inst_cellmath__47_0_in4), .D(inst_cellmath__47_0_in0));
NOR2XL inst_cellmath__47_0_I5 (.Y(inst_cellmath__47_0_out0), .A(N12), .B(inst_cellmath__47_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__53_U_bdw2876250654_bdw (
	inst_cellmath__53_U_out0,
	inst_cellmath__53_U_in0,
	inst_cellmath__53_U_in1,
	inst_cellmath__53_U_in2,
	inst_cellmath__53_U_in3,
	inst_cellmath__53_U_in4,
	inst_cellmath__53_U_in5
	); /* architecture "gate_level" */ 
output [22:22] inst_cellmath__53_U_out0;
input  inst_cellmath__53_U_in0,
	inst_cellmath__53_U_in1;
input [22:22] inst_cellmath__53_U_in2;
input  inst_cellmath__53_U_in3,
	inst_cellmath__53_U_in4;
input [46:46] inst_cellmath__53_U_in5;
wire N13,N17;
NOR2XL inst_cellmath__53_U_I1 (.Y(N13), .A(inst_cellmath__53_U_in4), .B(inst_cellmath__53_U_in1));
MXI2XL inst_cellmath__53_U_I6 (.Y(N17), .A(inst_cellmath__53_U_in5[46]), .B(inst_cellmath__53_U_in2[22]), .S0(inst_cellmath__53_U_in3));
MXI2XL inst_cellmath__53_U_I7 (.Y(inst_cellmath__53_U_out0[22]), .A(N17), .B(N13), .S0(inst_cellmath__53_U_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2876250654_bdw (
	inst_cellmath__53_M_out0,
	inst_cellmath__53_M_in0,
	inst_cellmath__53_M_in1,
	inst_cellmath__53_M_in2,
	inst_cellmath__53_M_in3,
	inst_cellmath__53_M_in4,
	inst_cellmath__53_M_in5,
	inst_cellmath__53_M_in6,
	inst_cellmath__53_M_in7,
	inst_cellmath__53_M_in8,
	inst_cellmath__53_M_in9
	); /* architecture "gate_level" */ 
output [21:0] inst_cellmath__53_M_out0;
input  inst_cellmath__53_M_in0,
	inst_cellmath__53_M_in1;
input [21:0] inst_cellmath__53_M_in2;
input  inst_cellmath__53_M_in3,
	inst_cellmath__53_M_in4;
input [45:24] inst_cellmath__53_M_in5;
input  inst_cellmath__53_M_in6,
	inst_cellmath__53_M_in7;
input [21:0] inst_cellmath__53_M_in8,
	inst_cellmath__53_M_in9;
wire N135,N137,N142,N144,N146,N148,N150 
	,N152,N154,N156,N158,N160,N162,N164,N166 
	,N168,N170,N172,N174,N176,N178,N180,N182 
	,N184,N236,N238,N240,N242,N244,N246,N248 
	,N250,N252,N254,N256,N258,N260,N262,N264 
	,N266,N268,N270,N272,N274,N276,N278,N281 
	,N285,N289,N293,N297,N301,N305,N309,N313 
	,N317,N321,N325,N329,N333,N337,N341,N345 
	,N349,N353,N357,N361,N365,N368,N370,N372 
	,N538,N547,N548;
INVXL inst_cellmath__53_M_I182 (.Y(N538), .A(inst_cellmath__53_M_in0));
NOR2XL inst_cellmath__53_M_I7 (.Y(N368), .A(inst_cellmath__53_M_in4), .B(N538));
NAND3BXL inst_cellmath__53_M_I429 (.Y(N135), .AN(inst_cellmath__53_M_in7), .B(inst_cellmath__53_M_in6), .C(inst_cellmath__53_M_in4));
NOR2XL inst_cellmath__53_M_I11 (.Y(N370), .A(N135), .B(N538));
NAND2XL inst_cellmath__53_M_I12 (.Y(N137), .A(inst_cellmath__53_M_in7), .B(inst_cellmath__53_M_in4));
NOR2XL inst_cellmath__53_M_I13 (.Y(N372), .A(N137), .B(N538));
NOR2BX1 inst_cellmath__53_M_I200 (.Y(N547), .AN(N538), .B(inst_cellmath__53_M_in3));
AND2XL inst_cellmath__53_M_I201 (.Y(N548), .A(inst_cellmath__53_M_in3), .B(N538));
AOI22XL inst_cellmath__53_M_I17 (.Y(N142), .A0(inst_cellmath__53_M_in2[0]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[24]));
AOI22XL inst_cellmath__53_M_I18 (.Y(N144), .A0(inst_cellmath__53_M_in2[1]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[25]));
AOI22XL inst_cellmath__53_M_I19 (.Y(N146), .A0(inst_cellmath__53_M_in2[2]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[26]));
AOI22XL inst_cellmath__53_M_I20 (.Y(N148), .A0(inst_cellmath__53_M_in2[3]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[27]));
AOI22XL inst_cellmath__53_M_I21 (.Y(N150), .A0(inst_cellmath__53_M_in2[4]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[28]));
AOI22XL inst_cellmath__53_M_I22 (.Y(N152), .A0(inst_cellmath__53_M_in2[5]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[29]));
AOI22XL inst_cellmath__53_M_I23 (.Y(N154), .A0(inst_cellmath__53_M_in2[6]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[30]));
AOI22XL inst_cellmath__53_M_I24 (.Y(N156), .A0(inst_cellmath__53_M_in2[7]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[31]));
AOI22XL inst_cellmath__53_M_I25 (.Y(N158), .A0(inst_cellmath__53_M_in2[8]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[32]));
AOI22XL inst_cellmath__53_M_I26 (.Y(N160), .A0(inst_cellmath__53_M_in2[9]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[33]));
AOI22XL inst_cellmath__53_M_I27 (.Y(N162), .A0(inst_cellmath__53_M_in2[10]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[34]));
AOI22XL inst_cellmath__53_M_I28 (.Y(N164), .A0(inst_cellmath__53_M_in2[11]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[35]));
AOI22XL inst_cellmath__53_M_I29 (.Y(N166), .A0(inst_cellmath__53_M_in2[12]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[36]));
AOI22XL inst_cellmath__53_M_I30 (.Y(N168), .A0(inst_cellmath__53_M_in2[13]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[37]));
AOI22XL inst_cellmath__53_M_I31 (.Y(N170), .A0(inst_cellmath__53_M_in2[14]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[38]));
AOI22XL inst_cellmath__53_M_I32 (.Y(N172), .A0(inst_cellmath__53_M_in2[15]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[39]));
AOI22XL inst_cellmath__53_M_I33 (.Y(N174), .A0(inst_cellmath__53_M_in2[16]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[40]));
AOI22XL inst_cellmath__53_M_I34 (.Y(N176), .A0(inst_cellmath__53_M_in2[17]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[41]));
AOI22XL inst_cellmath__53_M_I35 (.Y(N178), .A0(inst_cellmath__53_M_in2[18]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[42]));
AOI22XL inst_cellmath__53_M_I36 (.Y(N180), .A0(inst_cellmath__53_M_in2[19]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[43]));
AOI22XL inst_cellmath__53_M_I37 (.Y(N182), .A0(inst_cellmath__53_M_in2[20]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[44]));
AOI22XL inst_cellmath__53_M_I38 (.Y(N184), .A0(inst_cellmath__53_M_in2[21]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[45]));
AOI22XL inst_cellmath__53_M_I42 (.Y(N281), .A0(inst_cellmath__53_M_in8[0]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I43 (.Y(N285), .A0(inst_cellmath__53_M_in8[1]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I44 (.Y(N289), .A0(inst_cellmath__53_M_in8[2]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I45 (.Y(N293), .A0(inst_cellmath__53_M_in8[3]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I46 (.Y(N297), .A0(inst_cellmath__53_M_in8[4]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I47 (.Y(N301), .A0(inst_cellmath__53_M_in8[5]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I48 (.Y(N305), .A0(inst_cellmath__53_M_in8[6]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I49 (.Y(N309), .A0(inst_cellmath__53_M_in8[7]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I50 (.Y(N313), .A0(inst_cellmath__53_M_in8[8]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I51 (.Y(N317), .A0(inst_cellmath__53_M_in8[9]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I52 (.Y(N321), .A0(inst_cellmath__53_M_in8[10]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I53 (.Y(N325), .A0(inst_cellmath__53_M_in8[11]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I54 (.Y(N329), .A0(inst_cellmath__53_M_in8[12]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I55 (.Y(N333), .A0(inst_cellmath__53_M_in8[13]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I56 (.Y(N337), .A0(inst_cellmath__53_M_in8[14]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I57 (.Y(N341), .A0(inst_cellmath__53_M_in8[15]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I58 (.Y(N345), .A0(inst_cellmath__53_M_in8[16]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I59 (.Y(N349), .A0(inst_cellmath__53_M_in8[17]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I60 (.Y(N353), .A0(inst_cellmath__53_M_in8[18]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I61 (.Y(N357), .A0(inst_cellmath__53_M_in8[19]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I62 (.Y(N361), .A0(inst_cellmath__53_M_in8[20]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I63 (.Y(N365), .A0(inst_cellmath__53_M_in8[21]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
NAND2XL inst_cellmath__53_M_I67 (.Y(N236), .A(N372), .B(inst_cellmath__53_M_in9[0]));
NAND2XL inst_cellmath__53_M_I68 (.Y(N238), .A(N372), .B(inst_cellmath__53_M_in9[1]));
NAND2XL inst_cellmath__53_M_I69 (.Y(N240), .A(N372), .B(inst_cellmath__53_M_in9[2]));
NAND2XL inst_cellmath__53_M_I70 (.Y(N242), .A(N372), .B(inst_cellmath__53_M_in9[3]));
NAND2XL inst_cellmath__53_M_I71 (.Y(N244), .A(N372), .B(inst_cellmath__53_M_in9[4]));
NAND2XL inst_cellmath__53_M_I72 (.Y(N246), .A(N372), .B(inst_cellmath__53_M_in9[5]));
NAND2XL inst_cellmath__53_M_I73 (.Y(N248), .A(N372), .B(inst_cellmath__53_M_in9[6]));
NAND2XL inst_cellmath__53_M_I74 (.Y(N250), .A(N372), .B(inst_cellmath__53_M_in9[7]));
NAND2XL inst_cellmath__53_M_I75 (.Y(N252), .A(N372), .B(inst_cellmath__53_M_in9[8]));
NAND2XL inst_cellmath__53_M_I76 (.Y(N254), .A(N372), .B(inst_cellmath__53_M_in9[9]));
NAND2XL inst_cellmath__53_M_I77 (.Y(N256), .A(N372), .B(inst_cellmath__53_M_in9[10]));
NAND2XL inst_cellmath__53_M_I78 (.Y(N258), .A(N372), .B(inst_cellmath__53_M_in9[11]));
NAND2XL inst_cellmath__53_M_I79 (.Y(N260), .A(N372), .B(inst_cellmath__53_M_in9[12]));
NAND2XL inst_cellmath__53_M_I80 (.Y(N262), .A(N372), .B(inst_cellmath__53_M_in9[13]));
NAND2XL inst_cellmath__53_M_I81 (.Y(N264), .A(N372), .B(inst_cellmath__53_M_in9[14]));
NAND2XL inst_cellmath__53_M_I82 (.Y(N266), .A(N372), .B(inst_cellmath__53_M_in9[15]));
NAND2XL inst_cellmath__53_M_I83 (.Y(N268), .A(N372), .B(inst_cellmath__53_M_in9[16]));
NAND2XL inst_cellmath__53_M_I84 (.Y(N270), .A(N372), .B(inst_cellmath__53_M_in9[17]));
NAND2XL inst_cellmath__53_M_I85 (.Y(N272), .A(N372), .B(inst_cellmath__53_M_in9[18]));
NAND2XL inst_cellmath__53_M_I86 (.Y(N274), .A(N372), .B(inst_cellmath__53_M_in9[19]));
NAND2XL inst_cellmath__53_M_I87 (.Y(N276), .A(N372), .B(inst_cellmath__53_M_in9[20]));
NAND2XL inst_cellmath__53_M_I88 (.Y(N278), .A(N372), .B(inst_cellmath__53_M_in9[21]));
NAND3XL inst_cellmath__53_M_I202 (.Y(inst_cellmath__53_M_out0[0]), .A(N236), .B(N142), .C(N281));
NAND3XL inst_cellmath__53_M_I203 (.Y(inst_cellmath__53_M_out0[1]), .A(N238), .B(N144), .C(N285));
NAND3XL inst_cellmath__53_M_I204 (.Y(inst_cellmath__53_M_out0[2]), .A(N240), .B(N146), .C(N289));
NAND3XL inst_cellmath__53_M_I205 (.Y(inst_cellmath__53_M_out0[3]), .A(N242), .B(N148), .C(N293));
NAND3XL inst_cellmath__53_M_I206 (.Y(inst_cellmath__53_M_out0[4]), .A(N244), .B(N150), .C(N297));
NAND3XL inst_cellmath__53_M_I207 (.Y(inst_cellmath__53_M_out0[5]), .A(N246), .B(N152), .C(N301));
NAND3XL inst_cellmath__53_M_I208 (.Y(inst_cellmath__53_M_out0[6]), .A(N248), .B(N154), .C(N305));
NAND3XL inst_cellmath__53_M_I209 (.Y(inst_cellmath__53_M_out0[7]), .A(N250), .B(N156), .C(N309));
NAND3XL inst_cellmath__53_M_I210 (.Y(inst_cellmath__53_M_out0[8]), .A(N252), .B(N158), .C(N313));
NAND3XL inst_cellmath__53_M_I211 (.Y(inst_cellmath__53_M_out0[9]), .A(N254), .B(N160), .C(N317));
NAND3XL inst_cellmath__53_M_I212 (.Y(inst_cellmath__53_M_out0[10]), .A(N256), .B(N162), .C(N321));
NAND3XL inst_cellmath__53_M_I213 (.Y(inst_cellmath__53_M_out0[11]), .A(N258), .B(N164), .C(N325));
NAND3XL inst_cellmath__53_M_I214 (.Y(inst_cellmath__53_M_out0[12]), .A(N260), .B(N166), .C(N329));
NAND3XL inst_cellmath__53_M_I215 (.Y(inst_cellmath__53_M_out0[13]), .A(N262), .B(N168), .C(N333));
NAND3XL inst_cellmath__53_M_I216 (.Y(inst_cellmath__53_M_out0[14]), .A(N264), .B(N170), .C(N337));
NAND3XL inst_cellmath__53_M_I217 (.Y(inst_cellmath__53_M_out0[15]), .A(N266), .B(N172), .C(N341));
NAND3XL inst_cellmath__53_M_I218 (.Y(inst_cellmath__53_M_out0[16]), .A(N268), .B(N174), .C(N345));
NAND3XL inst_cellmath__53_M_I219 (.Y(inst_cellmath__53_M_out0[17]), .A(N270), .B(N176), .C(N349));
NAND3XL inst_cellmath__53_M_I220 (.Y(inst_cellmath__53_M_out0[18]), .A(N272), .B(N178), .C(N353));
NAND3XL inst_cellmath__53_M_I221 (.Y(inst_cellmath__53_M_out0[19]), .A(N274), .B(N180), .C(N357));
NAND3XL inst_cellmath__53_M_I222 (.Y(inst_cellmath__53_M_out0[20]), .A(N276), .B(N182), .C(N361));
NAND3XL inst_cellmath__53_M_I223 (.Y(inst_cellmath__53_M_out0[21]), .A(N278), .B(N184), .C(N365));
endmodule

/* CADENCE  ubH2TQzarhA= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




module float_div_cynw_cm_float_mul_ieee_E8_M23_3_0( a_sign, a_exp, a_man, b_sign, b_exp, b_man, rm, x, aclk, astall );
input a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire[31:0] x_wire;
input aclk;
input astall;
cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2876250654_bdw cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw3828364039_bdw_inst( .a_sign(a_sign), .a_exp(a_exp), .a_man(a_man), .b_sign(b_sign), .b_exp(b_exp), .b_man(b_man), .rm(rm), .x(x_wire));
reg [31:0] x_reg_0;
/* $A : movable_reg */
always @(posedge aclk) begin
    if ( !astall) x_reg_0 <= x_wire;
end
/* $A : movable_reg = reset */
assign x = x_reg_0;
endmodule


