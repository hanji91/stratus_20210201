/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:04 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_5 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51;
wire [24:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2695,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2696,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2720,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2865,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7520,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7646,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7980,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795;
wire N5677,N5682,N5687,N5692,N5697,N5702,N5707 
	,N5712,N5717,N11884,N11888,N11890,N12051,N12056,N12061 
	,N12066,N12071,N12076,N12164,N12168,N12170,N12229,N12234 
	,N12239,N12244,N12249,N12254,N12259,N12266,N12274,N12291 
	,N12295,N12309,N12317,N12325,N12333,N12349,N12365,N12416 
	,N12418,N12420,N12445,N12449,N12511,N12513,N12546,N12581 
	,N12587,N12589,N12622,N12628,N12663,N12704,N12724,N12726 
	,N12728,N12769,N12777,N12781,N12822,N12881,N12895,N12945 
	,N12967,N12975,N12977,N12979,N13040,N13048,N13060,N13066 
	,N13068,N13070,N13129,N13145,N13153,N13155,N13157,N13215 
	,N13223,N13235,N13241,N13243,N13245,N13254,N13261,N13263 
	,N13319,N13364,N13366,N13432,N13455,N13465,N13470,N13476 
	,N13478,N13494,N13496,N13498,N13610,N13616,N13618,N13624 
	,N13626,N13628,N13706,N13712,N13720,N13727,N13735,N13745 
	,N13751,N13753,N13755,N13759,N13761,N13767,N13769,N13771 
	,N13780,N13782,N13784,N13849,N13859,N13867,N13869,N13883 
	,N13885,N13889,N13907,N13917,N13925,N13931,N13933,N13935 
	,N13944,N13946,N13948,N14002,N14006,N14014,N14018,N14024 
	,N14030,N14038,N14040,N14060,N14071,N14073,N14075,N14079 
	,N14081,N14083,N14087,N14089,N14091,N14158,N14160,N14166 
	,N14168,N14174,N14178,N14182,N14184,N14186,N14202,N14204 
	,N14206,N14209,N14214,N14230,N14232,N14234,N14260,N14278 
	,N14284,N14286,N14288,N14292,N14294,N14296,N14301,N14316 
	,N14318,N14320,N14324,N14326,N14328,N14339,N14370,N14374 
	,N14376,N14378,N14382,N14384,N14386,N14390,N14392,N14394 
	,N14398,N14400,N14402,N14406,N14408,N14419,N14421,N14423 
	,N14435,N14441,N14443,N14454,N14456,N14465,N14469,N14471 
	,N14473,N14479,N14481,N14483,N14487,N14489,N14491,N14494 
	,N14505,N14507,N14509,N14515,N14517,N14519,N14526,N14535 
	,N14543,N14551,N14556,N14562,N15230,N15238,N15245,N15271 
	,N15281,N15285,N15287,N15289,N15293,N15832,N15834,N15845 
	,N15848,N15849,N15851,N15853,N15854,N15856,N15858,N15860 
	,N15861,N15863,N15865,N15867,N15869,N15870,N15871,N15873 
	,N15875,N15878,N15881,N15883,N15885,N15886,N15888,N15894 
	,N15929,N15933,N15934,N15935,N15936,N15939,N15940,N15942 
	,N15944,N15947,N15949,N15952,N15957,N15959,N15963,N15993 
	,N15996,N15997,N16001,N16003,N16005,N16008,N16010,N16012 
	,N16014,N16016,N16017,N16019,N16020,N16022,N16025,N16027 
	,N16029,N16030,N16032,N16034,N16038,N16039,N16040,N16042 
	,N16075,N16079,N16080,N16082,N16084,N16085,N16087,N16089 
	,N16091,N16093,N16095,N16099,N16101,N16102,N16104,N16105 
	,N16107,N16108,N16111,N16113,N16115,N16116,N16119,N16120 
	,N16121,N16123,N16126,N16128,N16162,N16165,N16167,N16168 
	,N16169,N16171,N16173,N16185,N16186,N16190,N16193,N16194 
	,N16197,N16199,N16201,N16203;
EDFFHQX1 x_reg_L1_22__retimed_I8255 (.Q(N15293), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I8254 (.Q(x[13]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8253 (.Q(N15289), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8252 (.Q(N15287), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8251 (.Q(N15285), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8250 (.Q(N15281), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8246 (.Q(N15271), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2803), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8235 (.Q(N15245), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8232 (.Q(N15238), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I8229 (.Q(N15230), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7935 (.Q(N14519), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7934 (.Q(N14517), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7933 (.Q(N14515), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7932 (.Q(N14509), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7931 (.Q(N14507), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7930 (.Q(N14505), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7926 (.Q(N14494), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7925 (.Q(N14491), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7924 (.Q(N14489), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7923 (.Q(N14487), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7922 (.Q(N14483), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7921 (.Q(N14481), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7920 (.Q(N14479), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7919 (.Q(N14473), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7918 (.Q(N14471), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7917 (.Q(N14469), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7916 (.Q(N14465), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7912 (.Q(N14456), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7911 (.Q(N14454), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7907 (.Q(N14443), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7906 (.Q(N14441), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7905 (.Q(N14435), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7904 (.Q(N14423), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7903 (.Q(N14421), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7902 (.Q(N14419), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7898 (.Q(N14408), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7897 (.Q(N14406), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7896 (.Q(N14402), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7895 (.Q(N14400), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7894 (.Q(N14398), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7893 (.Q(N14394), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7892 (.Q(N14392), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7891 (.Q(N14390), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7890 (.Q(N14386), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7889 (.Q(N14384), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7888 (.Q(N14382), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7887 (.Q(N14378), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7886 (.Q(N14376), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7885 (.Q(N14374), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7884 (.Q(N14370), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7871 (.Q(N14339), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7868 (.Q(N14328), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7867 (.Q(N14326), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7866 (.Q(N14324), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7865 (.Q(N14320), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7864 (.Q(N14318), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7863 (.Q(N14316), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7861 (.Q(N14301), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2588), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7859 (.Q(N14296), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7858 (.Q(N14294), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7857 (.Q(N14292), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7856 (.Q(N14288), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7855 (.Q(N14286), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7854 (.Q(N14284), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7852 (.Q(N14278), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7845 (.Q(N14260), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7836 (.Q(N14234), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7835 (.Q(N14232), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7834 (.Q(N14230), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7828 (.Q(N14214), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7826 (.Q(N14209), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7825 (.Q(N14206), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7824 (.Q(N14204), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7823 (.Q(N14202), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7821 (.Q(N14186), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7820 (.Q(N14184), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7819 (.Q(N14182), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7818 (.Q(N14178), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7816 (.Q(N14174), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7814 (.Q(N14168), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7813 (.Q(N14166), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7811 (.Q(N14160), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7810 (.Q(N14158), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7785 (.Q(N14091), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7784 (.Q(N14089), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7783 (.Q(N14087), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7782 (.Q(N14083), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7781 (.Q(N14081), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7780 (.Q(N14079), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7779 (.Q(N14075), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7778 (.Q(N14073), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7777 (.Q(N14071), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7773 (.Q(N14060), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7765 (.Q(N14040), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7764 (.Q(N14038), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7761 (.Q(N14030), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7759 (.Q(N14024), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7757 (.Q(N14018), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7755 (.Q(N14014), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7752 (.Q(N14006), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7751 (.Q(N14002), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7731 (.Q(N13948), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7730 (.Q(N13946), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7729 (.Q(N13944), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7726 (.Q(N13935), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7725 (.Q(N13933), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7724 (.Q(N13931), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7722 (.Q(N13925), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7719 (.Q(N13917), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7715 (.Q(N13907), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7708 (.Q(N13889), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7707 (.Q(N13885), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7706 (.Q(N13883), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7701 (.Q(N13869), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7700 (.Q(N13867), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7697 (.Q(N13859), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7693 (.Q(N13849), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7669 (.Q(N13784), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7668 (.Q(N13782), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7667 (.Q(N13780), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7664 (.Q(N13771), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7663 (.Q(N13769), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7662 (.Q(N13767), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7660 (.Q(N13761), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7659 (.Q(N13759), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7658 (.Q(N13755), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7657 (.Q(N13753), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7656 (.Q(N13751), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7654 (.Q(N13745), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7650 (.Q(N13735), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7647 (.Q(N13727), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7645 (.Q(N13720), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7642 (.Q(N13712), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7640 (.Q(N13706), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7611 (.Q(N13628), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7610 (.Q(N13626), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7609 (.Q(N13624), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7607 (.Q(N13618), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7606 (.Q(N13616), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7604 (.Q(N13610), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7562 (.Q(N13498), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7561 (.Q(N13496), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7560 (.Q(N13494), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7554 (.Q(N13478), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7553 (.Q(N13476), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7551 (.Q(N13470), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7549 (.Q(N13465), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7545 (.Q(N13455), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7536 (.Q(N13432), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7512 (.Q(N13366), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7511 (.Q(N13364), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7494 (.Q(N13319), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I7474 (.Q(N13263), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I7473 (.Q(N13261), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7470 (.Q(N13254), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7467 (.Q(N13245), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7466 (.Q(N13243), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7465 (.Q(N13241), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7463 (.Q(N13235), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7458 (.Q(N13223), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7455 (.Q(N13215), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7434 (.Q(N13157), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7433 (.Q(N13155), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7432 (.Q(N13153), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7429 (.Q(N13145), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7423 (.Q(N13129), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7402 (.Q(N13070), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7401 (.Q(N13068), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7400 (.Q(N13066), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7398 (.Q(N13060), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7393 (.Q(N13048), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7390 (.Q(N13040), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7369 (.Q(N12979), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7368 (.Q(N12977), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7367 (.Q(N12975), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7364 (.Q(N12967), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7356 (.Q(N12945), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7338 (.Q(N12895), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7333 (.Q(N12881), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7312 (.Q(N12822), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7298 (.Q(N12781), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7296 (.Q(N12777), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7293 (.Q(N12769), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7279 (.Q(N12728), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7278 (.Q(N12726), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7277 (.Q(N12724), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7270 (.Q(N12704), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7256 (.Q(N12663), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7244 (.Q(N12628), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7242 (.Q(N12622), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7231 (.Q(N12589), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7230 (.Q(N12587), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7228 (.Q(N12581), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7216 (.Q(N12546), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7205 (.Q(N12513), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7204 (.Q(N12511), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7183 (.Q(N12449), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7181 (.Q(N12445), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7173 (.Q(N12420), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7172 (.Q(N12418), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7171 (.Q(N12416), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7153 (.Q(N12365), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7147 (.Q(N12349), .D(N12325), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7141 (.Q(N12333), .D(N12309), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7138 (.Q(N12325), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7135 (.Q(N12317), .D(N12295), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7132 (.Q(N12309), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7127 (.Q(N12295), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7126 (.Q(N12291), .D(N12274), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7120 (.Q(N12274), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_14__retimed_I7117 (.Q(N12266), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_16__retimed_I7114 (.Q(N12259), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_17__retimed_I7112 (.Q(N12254), .D(N12076), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_18__retimed_I7110 (.Q(N12249), .D(N12071), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_19__retimed_I7108 (.Q(N12244), .D(N12066), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_20__retimed_I7106 (.Q(N12239), .D(N12061), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I7104 (.Q(N12234), .D(N12056), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7102 (.Q(N12229), .D(N12051), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7077 (.Q(N12170), .D(N11890), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7076 (.Q(N12168), .D(N11888), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I7074 (.Q(N12164), .D(N11884), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_17__retimed_I7039 (.Q(N12076), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_18__retimed_I7037 (.Q(N12071), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_19__retimed_I7035 (.Q(N12066), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_20__retimed_I7033 (.Q(N12061), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I7031 (.Q(N12056), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I7029 (.Q(N12051), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I6960 (.Q(N11890), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I6959 (.Q(N11888), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I6957 (.Q(N11884), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795), .E(bdw_enable), .CK(aclk));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_5_I0 (.Y(bdw_enable), .A(astall));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353), .A(a_exp[7]), .B(a_exp[0]));
AND4XL float_div_cynw_cm_float_rcp_E8_M23_5_I2 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL float_div_cynw_cm_float_rcp_E8_M23_5_I3 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743), .A(a_exp[6]), .B(a_exp[5]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I4 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I5 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376), .A(a_man[10]), .B(a_man[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I6 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395), .A(a_man[6]), .B(a_man[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I7 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384), .A(a_man[8]), .B(a_man[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404), .A(a_man[4]), .B(a_man[3]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_5_I9 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_5_I10 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_5_I11 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I12 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .A(a_man[18]), .B(a_man[17]));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_5_I13 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_5_I14 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B(a_man[16]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408), .D(a_man[15]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I15 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I16 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_5_I17 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I18 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I19 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I20 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I21 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_5_I22 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I23 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I24 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]), .A(a_exp[1]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I25 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0]), .A(a_exp[0]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I26 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I27 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I28 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]), .A(a_exp[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I29 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]), .A(a_exp[3]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I30 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457), .A(a_exp[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I31 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I32 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]), .A(a_exp[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I33 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I34 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451), .A(a_exp[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I35 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_5_I36 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I37 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I38 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]), .A(a_exp[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I39 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]), .A(a_exp[7]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I40 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444), .A(a_exp[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I41 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I42 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I43 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]), .A(a_exp[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I44 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_5_I45 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I46 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_5_I47 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8]));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I48 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_5_I49 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_5_I50 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I51 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I52 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I53 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I54 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A(a_man[21]));
CLKINVX4 float_div_cynw_cm_float_rcp_E8_M23_5_I55 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I56 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I57 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310), .B(a_man[20]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_5_I58 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A(a_man[20]));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_5_I59 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A(a_man[18]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I60 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .A(a_man[16]), .B(a_man[17]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I61 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I62 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I63 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I64 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071), .B1(a_man[21]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I65 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .A(a_man[17]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I66 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .A(a_man[16]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I67 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I68 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I69 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I70 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I71 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I72 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I73 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I74 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I75 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I76 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .A(a_man[17]), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I77 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I78 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I79 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I80 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I81 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I82 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .A(a_man[17]), .B(a_man[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I83 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_5_I84 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .A1N(a_man[19]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I85 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I86 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I87 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I88 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I89 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I90 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I91 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I92 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I93 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I94 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I95 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I96 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I97 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I98 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I99 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809), .B1(a_man[21]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022), .B0(a_man[19]), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054), .A(a_man[19]), .B(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I109 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I110 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I111 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_5_I113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[18]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213), .B1(a_man[22]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B1(a_man[19]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .A(a_man[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_5_I142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .A0(a_man[16]), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I145 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I161 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I162 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I166 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783), .A(1'B1), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I167 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I168 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I169 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I170 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .A(a_man[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I172 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I173 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400), .B1(a_man[20]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_5_I201 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589), .A1N(a_man[21]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I203 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .A(a_man[14]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I207 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]));
INVX1 gena_A_I8572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .A(a_man[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I213 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I214 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I215 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I216 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I217 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I221 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603), .B0(a_man[18]), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637), .A(a_man[12]));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_5_I242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848), .B(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I253 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888), .A(a_man[11]));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_5_I256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I258 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[18]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I259 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I260 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I269 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I271 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I272 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I273 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I274 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I275 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I276 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I289 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I290 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I291 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I293 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I300 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .A(a_man[10]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I302 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I303 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I304 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I305 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I310 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I314 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I315 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I318 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I319 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I323 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I324 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I325 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I326 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I327 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I328 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I329 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809), .A(N12418), .B(N12416), .CI(N12420));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006), .A(N12365), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I333 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I334 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I340 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I345 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I346 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I347 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I348 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I349 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I350 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I351 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I353 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I354 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747), .A(a_man[9]));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_5_I355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I371 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I372 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I373 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I377 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I378 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648), .A(a_man[8]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I382 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I384 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I385 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I387 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I388 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I389 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I390 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I391 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572), .A(N12511), .B(N12513));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I392 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892), .B(N12445), .CI(N12449));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I393 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I398 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I404 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I409 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I417 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8542 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .A(a_man[7]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I423 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I424 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I428 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I429 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I432 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I433 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I438 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I439 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I440 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I443 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I444 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I445 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I446 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I447 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I448 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I449 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I450 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I456 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I458 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I459 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I460 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I461 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I462 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I463 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I464 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B0(a_man[18]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I469 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I471 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I472 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I473 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I474 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I475 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I476 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .A(a_man[6]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I481 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I485 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I486 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I487 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I488 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I489 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I490 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I491 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I494 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I495 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I496 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I497 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I498 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I499 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I500 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I501 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I502 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I503 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I504 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I505 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888), .A(N12587), .B(N12589));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I506 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674), .A(N12546), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I507 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I508 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I509 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I510 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I517 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I518 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I520 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I522 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I523 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I524 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I525 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B(a_man[18]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I526 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I527 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I528 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I529 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I530 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I531 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I532 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I533 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I534 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I535 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I536 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I537 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I540 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I541 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I542 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I543 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I544 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I547 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698), .A(a_man[5]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I548 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I549 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I552 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I553 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I554 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I555 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I557 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I558 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I559 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I560 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I561 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I563 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I564 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I565 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I566 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I567 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I568 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I571 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I573 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I575 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I576 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I577 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I578 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I579 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]), .A(N12726), .B(N12724), .CI(N12728));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I580 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965), .A(N12628), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I581 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776), .A(N12581), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I582 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I583 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I584 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I585 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I587 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I588 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I589 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I592 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I593 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I594 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I596 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I598 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I600 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I601 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I602 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I605 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I606 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I607 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I608 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I609 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I610 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I611 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I612 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I613 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I614 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I615 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I616 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I617 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I618 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I619 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631), .A(a_man[4]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .A(a_man[3]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I626 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I627 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I629 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I630 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I632 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I633 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I636 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I637 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I638 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I639 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I640 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I641 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I642 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I643 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I644 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I645 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I646 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I647 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I648 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I649 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I650 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I651 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I652 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I653 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I654 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I655 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I656 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I657 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I661 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I666 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I667 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I669 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I671 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I672 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I675 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I676 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I677 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I679 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I680 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I681 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I682 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I686 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I687 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I688 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I690 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I691 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I692 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I693 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I694 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530), .A(N15287), .B(N15285), .CI(N15289));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I695 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I696 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854), .B(N12777), .CI(N12781));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I697 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I698 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876), .A(N12622), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I699 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I700 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I701 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I702 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I704 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I705 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I706 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I707 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I708 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I709 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I710 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I711 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I712 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I713 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I714 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I715 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I719 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I721 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I723 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I724 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I725 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I726 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I727 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I728 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I729 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I730 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I731 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I733 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .A(a_man[2]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I734 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .A(a_man[0]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I735 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .A(a_man[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I736 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I737 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I738 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I739 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I740 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I741 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I742 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I746 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I747 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I748 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I749 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105), .A(N12977), .B(N12975), .CI(N12979));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I750 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294), .B(N12769), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I751 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I752 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982), .A(N12663), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I753 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I754 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I755 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I756 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I757 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467));
INVXL gena_A_I8573 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I765 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2853), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I766 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2831), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I767 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I768 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I769 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I770 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2706), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2638), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I773 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I774 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I775 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I777 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2784), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8544 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2748), .S(N15860), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I778 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2748), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2784), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2638));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I781 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I782 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I785 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I786 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I787 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I789 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8545 (.CO(N15894), .S(N15886), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8546 (.CO(N15865), .S(N15853), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8547 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889), .S(N15878), .A(N15860), .B(N15894), .CI(N15865));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I792 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I793 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I794 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I795 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I796 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I798 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I799 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I800 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I801 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I805 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I806 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I807 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I808 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I809 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I812 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I813 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I814 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I815 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I816 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I817 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I818 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I819 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I820 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I821 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I822 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I823 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I825 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I826 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2865), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I827 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I828 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I829 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I831 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I832 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I833 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I834 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I835 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I837 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I838 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I839 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I840 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I841 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8597 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2880), .S(N15996), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I843 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2683), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2880));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I844 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I845 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I846 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I847 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I848 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I850 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I852 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I853 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I854 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I855 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8598 (.CO(N16030), .S(N16016), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8599 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2695), .S(N16042), .A(N16030), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I857 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2695), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2865), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2683));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I858 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I859 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I860 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I861 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I862 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8600 (.CO(N16022), .S(N16008), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8601 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841), .S(N16034), .A(N16022), .B(N15996), .CI(N16042));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I865 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I866 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I867 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I868 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I869 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I870 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I871 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I876 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I877 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I879 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I883 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I884 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I885 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I886 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I887 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8622 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702), .S(N16079), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8602 (.CO(N16014), .S(N16003), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8623 (.CO(N16115), .S(N16101), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8624 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846), .S(N16128), .A(N16115), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8605 (.CO(N16020), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872), .CI(N16003));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8625 (.CO(N16107), .S(N16095), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8626 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660), .S(N16120), .A(N16079), .B(N16107), .CI(N16128));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I891 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I892 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I893 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I894 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I898 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I899 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I900 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I903 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I904 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I905 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I906 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I909 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I910 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I911 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I912 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I913 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I914 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8636 (.CO(N16087), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I918 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I919 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I920 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_5_I921 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I922 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I923 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I924 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I925 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I926 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8627 (.CO(N16099), .S(N16089), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8628 (.CO(N16126), .S(N16113), .A(N16099), .B(N16101), .CI(N16095));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8629 (.Y(N16085), .A(N16126));
MXI2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8630 (.Y(N16121), .A(N16126), .B(N16085), .S0(N16120));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8631 (.CO(N16105), .S(N16093), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726), .CI(N16089));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8632 (.Y(N16116), .A(N16105));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8633 (.Y(N16123), .A(N16116), .B(N16113));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8634 (.Y(N16084), .A(N16116), .B(N16113));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8635 (.Y(N16075), .A(N16084));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I8637 (.Y(N16111), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8638 (.Y(N16082), .A0(N16093), .A1(N16087), .B0(N16111));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8639 (.Y(N16108), .A(N16087), .B(N16093));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8640 (.Y(N16091), .A(N16108), .B(N16082));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8641 (.Y(N16080), .A(N16105), .B(N16113));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8642 (.Y(N16119), .A0(N16123), .A1(N16075), .B0(N16091));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8643 (.Y(N16104), .A(N16080), .B(N16119));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8644 (.Y(N16102), .A(N16126), .B(N16120));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I8645 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576), .A0(N16104), .A1(N16121), .B0(N16102));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8603 (.CO(N16039), .S(N16027), .A(N16016), .B(N16014), .CI(N16008));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652), .A(N16039), .B(N16034));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8606 (.Y(N16005), .A(N16020));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8607 (.Y(N16010), .A(N16005), .B(N16027));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8608 (.Y(N16029), .A(N16005), .B(N16027));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8609 (.Y(N16017), .A(N16029));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8610 (.Y(N16032), .A(N16020), .B(N16027));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8611 (.Y(N15993), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8612 (.Y(N16001), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8613 (.Y(N16012), .A(N15993), .B(N16001));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8614 (.Y(N16025), .A(N16020), .B(N16027));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8615 (.Y(N16040), .A0(N16010), .A1(N16017), .B0(N15993), .B1(N16001));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_5_I8616 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871), .A0(N16032), .A1(N16012), .B0(N16025));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8617 (.Y(N15997), .A(N16039), .B(N16034));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8618 (.Y(N16038), .A(N15997));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8619 (.Y(N16019), .A0(N16025), .A1(N16040), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749), .A(N16038), .B(N16019));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I939 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2720), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_5_I940 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2720));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_5_I942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I943 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8548 (.CO(N15858), .S(N15845), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8549 (.CO(N15883), .S(N15873), .A(N15858), .B(N15886), .CI(N15853));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852), .A(N15883), .B(N15878));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8551 (.CO(N15863), .S(N15851), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802), .CI(N15845));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8552 (.Y(N15861), .A(N15863));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8553 (.Y(N15867), .A(N15861), .B(N15873));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8554 (.Y(N15885), .A(N15861), .B(N15873));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8555 (.Y(N15875), .A(N15885));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710), .A(N15863), .B(N15873));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8557 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729), .B(N15851));
AO21X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8558 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8559 (.Y(N15856), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729), .B(N15851));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8560 (.Y(N15888), .A(N15856));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8561 (.Y(N15870), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_5_I8562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580), .B0(N15856));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8563 (.Y(N15854), .A(N15873));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8564 (.Y(N15881), .A(N15863), .B(N15873));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8565 (.Y(N15871), .A0(N15867), .A1(N15875), .B0(N15888), .B1(N15870));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_5_I8566 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627), .A0(N15854), .A1(N15861), .B0(N15871));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8567 (.Y(N15849), .A(N15883), .B(N15878));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8568 (.Y(N15869), .A(N15849));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I8569 (.Y(N15848), .A0(N15881), .A1(N15871), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703), .A(N15869), .B(N15848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I951 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2599), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778));
OR2XL gena_A_I8574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL gena_A_I8575 (.Y(N15963), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
INVXL gena_A_I8576 (.Y(N15934), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
OR2XL gena_A_I8577 (.Y(N15944), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
ADDFX1 gena_A_I8578 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809), .S(N15952), .A(N15963), .B(N15934), .CI(N15944));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I957 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2696), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809));
INVXL gena_A_I8518 (.Y(N15832), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2696));
XOR2XL gena_A_I8579 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809));
ADDFX1 gena_A_I8580 (.CO(N15947), .S(N15939), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2853), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2831), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2706));
INVXL gena_A_I8581 (.Y(N15929), .A(N15952));
NAND2XL gena_A_I8582 (.Y(N15933), .A(N15929), .B(N15947));
INVXL gena_A_I8583 (.Y(N15959), .A(N15947));
NAND2XL gena_A_I8584 (.Y(N15940), .A(N15952), .B(N15959));
XOR2XL gena_A_I8585 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625), .A(N15952), .B(N15947));
XOR2XL gena_A_I8586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813), .A(N15939), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849));
AO21XL gena_A_I8587 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2599));
NOR2XL gena_A_I8588 (.Y(N15942), .A(N15939), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849));
INVXL gena_A_I8589 (.Y(N15949), .A(N15942));
NAND2X1 gena_A_I8590 (.Y(N15935), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601));
AO21XL gena_A_I8591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601), .B0(N15942));
NOR2XL gena_A_I8592 (.Y(N15957), .A(N15952), .B(N15947));
AOI22X1 gena_A_I8593 (.Y(N15936), .A0(N15933), .A1(N15940), .B0(N15949), .B1(N15935));
AO21XL gena_A_I8594 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811), .A0(N15959), .A1(N15929), .B0(N15936));
OAI21XL gena_A_I8595 (.Y(N15834), .A0(N15957), .A1(N15936), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769));
NAND2XL gena_A_I8520 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2803), .A(N15832), .B(N15834));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_5_I959 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2588), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I960 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[24]), .A(N15271), .B(N14301));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I961 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[24]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I962 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24]), .A(N13060), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I963 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I964 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I965 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I966 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I967 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I968 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I969 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I970 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I971 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I972 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I973 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I974 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I975 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I979 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I980 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I982 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I983 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I984 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I985 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I986 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I987 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I989 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I990 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I991 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I992 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154), .A(N13235), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I993 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]), .A(N14406), .B(N14408));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_5_I994 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I995 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219), .A(N13060), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I996 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341), .A(N13235), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I997 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I998 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367), .A(N14435));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I999 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072), .A(N13060), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1000 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1001 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1002 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1003 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1004 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1005 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917), .A(a_man[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1006 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1007 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1008 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274), .A(N13470), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1009 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1010 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1011 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24]), .B(N12822), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1012 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1013 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1014 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1015 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1016 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1017 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1018 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1019 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1020 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1021 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1022 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1023 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1024 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1025 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1026 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1027 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1028 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1029 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1030 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1031 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1032 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1033 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1034 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1035 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1036 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1037 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1039 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1040 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1043 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1044 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1045 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1046 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1047 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1048 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1049 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1050 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1051 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1052 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1054 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1055 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1056 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1057 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1058 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1059 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1060 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1061 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1062 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1063 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1066 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1067 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1068 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1069 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1070 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1071 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1072 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1073 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1077 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1078 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1079 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1080 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332), .A(a_man[16]), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1081 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1082 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1085 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1086 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1087 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1088 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1089 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1090 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1091 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1092 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1095 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1096 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1097 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1098 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1099 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1105 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1108 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1109 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1110 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1111 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1136 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1140 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1145 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1146 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1151 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1155 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1159 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1160 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1161 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1162 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1163 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1164 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1165 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857), .A(N13155), .B(N13153), .CI(N13157));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1166 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1167 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169), .A(N13068), .B(N13066), .CI(N13070));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1168 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043), .B(N12967), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1169 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360), .B(N12895), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1170 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1171 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7459), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530), .B(N12704), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1172 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1173 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064), .B1(a_man[21]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1199 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1200 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1201 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1202 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1203 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1207 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1211 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1213 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1215 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1216 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1217 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1220 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1221 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1222 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1223 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1224 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031), .A(N13243), .B(N13241), .CI(N13245));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1225 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220), .B(N13048), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1226 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1227 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7937), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7565), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1228 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7937), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7459));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195), .A(N13235), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I1250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260), .A(N13060), .B(N15245));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127), .A(N13470), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1254 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318), .A(N13470), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387), .A(N13235), .B(N15245));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1258 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115), .A(N13060), .B(N15230));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1259 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1260 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1269 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401), .A(N13465), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1271 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1272 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1273 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7606), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7471), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23]), .B(N12881), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1274 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1275 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1276 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1289 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1290 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1291 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1293 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1300 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1302 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1303 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1304 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1305 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1310 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1314 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1315 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1318 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1319 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1323 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1324 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1325 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1326 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738), .A(N13496), .B(N13494), .CI(N13498));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1327 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833), .A(N13366), .B(N13364), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1328 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019), .B(N13145), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1329 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1333 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1334 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1340 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1345 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1346 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1347 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1348 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22]), .B(N12945), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1349 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7533), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7663), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7471), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1350 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7533), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7606), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7565));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1351 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1353 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1354 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378), .B1(a_man[20]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185), .A(N13745), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249), .A(N13465), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237), .A(N13235), .B(N15230));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1371 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196), .A(N13610), .B(N15281), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1372 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1373 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379), .A(N13745), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106), .A(N13465), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1377 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111), .B1(a_man[20]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1378 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1382 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1384 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1385 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1387 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1388 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1389 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310), .A(N13925), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1390 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1391 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1392 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1393 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1398 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1404 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1409 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1417 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1421 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1422 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1423 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1424 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1428 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1429 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1432 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1433 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1438 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1439 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1440 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1443 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1444 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1445 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1446 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1447 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511), .A(N13626), .B(N13624), .CI(N13628));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1448 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112), .A(N13478), .B(N13476), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1449 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299), .B(N13223), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1450 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1456 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1458 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1459 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1460 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1461 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1462 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1463 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1464 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1469 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1471 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21]), .B(N13040), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1472 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1473 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7663));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1474 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1475 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1476 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1481 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1485 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1486 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1487 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1488 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1489 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1490 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I1491 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1494 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1495 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1496 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1497 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1498 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037), .A(N13782), .B(N13780), .CI(N13784));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1499 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023), .A(N13618), .B(N13616), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1500 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1501 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1502 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1503 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1504 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1505 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1506 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[18]), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1507 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1508 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1509 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1510 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1517 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1518 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1520 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20]), .B(N13129), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1522 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1523 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1524 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1525 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1526 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1527 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1528 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1529 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1530 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1531 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1532 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1533 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1534 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1535 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1536 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1537 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1540 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1541 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1542 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1543 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094), .A(N15238), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1544 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355), .A(N13925), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081), .A(N13745), .B(N15245));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1547 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081), .CI(N13917));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1548 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283), .A(N13712), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1549 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1552 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326), .A(N13753), .B(N13751), .CI(N13755));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1553 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1554 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1555 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1557 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1558 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1559 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1560 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1561 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1563 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1564 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1565 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1566 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1567 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1568 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I1570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220), .A(N14060), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1571 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1573 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286), .A(N15238), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1575 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220), .B(N13889), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1576 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1577 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231), .A(N13745), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1578 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164), .A(N13925), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1579 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137), .A(N13720), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1580 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1581 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1582 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1583 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1584 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1585 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1586 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1587 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1588 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1589 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1592 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1593 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1594 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1596 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1598 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1600 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1601 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1602 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1605 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1606 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1607 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1608 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1609 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1610 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1611 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1612 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1613 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1614 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1615 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950), .A(N13946), .B(N13944), .CI(N13948));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1616 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415), .A(N13761), .B(N13759), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1617 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1618 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1619 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1626 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1627 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1629 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1630 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1632 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1633 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1636 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19]), .B(N13215), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1637 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270), .A(N13745), .B(N15230));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1638 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141), .A(N15238), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1639 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073), .A(N14060), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1640 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1641 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1642 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1643 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1644 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1645 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291), .A(N14081), .B(N14079), .CI(N14083));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1646 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364), .CI(N13706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1647 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1648 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262), .A(N14060), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1649 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1650 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1651 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1652 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1653 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1654 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1655 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1656 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1657 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1661 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197), .A(N14214), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1666 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269), .A(N14024), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1667 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1669 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1671 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123), .A(N14073), .B(N14071), .CI(N14075));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1672 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1675 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1676 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1677 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1679 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1680 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1681 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1682 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1686 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1687 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1688 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1690 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1691 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1692 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I1693 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1694 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129), .A(N14209), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1695 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1696 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1697 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1698 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1699 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080), .A(N13867), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129), .CI(N13869));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I1700 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342), .A(N14214), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1701 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1702 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1704 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1705 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246), .A(N13883), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342), .CI(N13885));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1706 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1707 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1708 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1709 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_5_I1710 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1711 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1712 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1713 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7969), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1714 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7980), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1715 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1719 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1721 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1723 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1724 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1725 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1726 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1727 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1728 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1729 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1730 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1731 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1733 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1734 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1735 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1736 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1737 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327), .A(N13769), .B(N13767), .CI(N13771));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1738 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1739 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1740 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1741 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1742 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1746 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1747 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1748 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1749 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1750 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1751 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1752 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1753 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1754 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1755 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1756 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1757 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18]), .B(N13319), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1758 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7771), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7450), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1759 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7771), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7980), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7969));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1760 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1762 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1763 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1764 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1765 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1766 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1767 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1768 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1769 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230), .A(N13933), .B(N13931), .CI(N13935));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1770 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1771 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1772 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1773 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1774 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1775 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1776 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1777 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1778 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1779 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1781 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1782 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1783 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1785 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1786 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17]), .B(N13432), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1787 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388), .A(N14214), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1789 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181), .A(N15238), .B(N15230));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1790 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388), .B(N14030), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I1791 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320), .A(N14209), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1792 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1793 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1794 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1795 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1796 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1798 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1799 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1800 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320), .B(N14014), .CI(N14018));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_5_I1801 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230), .A(N13859), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1802 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1803 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1804 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1805 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I1806 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174), .A(N14209), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1807 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086), .A(N14168), .B(N14166), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1808 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1809 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1810 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1811 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278), .A(N14204), .B(N14202), .CI(N14206));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1812 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354), .CI(N14002));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1813 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1814 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1815 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1816 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7649), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7520), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_5_I1817 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7984), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7561), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7520));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1818 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7984), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7649), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7450));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1819 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1820 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1821 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1822 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1823 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1825 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1826 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1827 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1828 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1829 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1831 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1832 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1833 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1834 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1835 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1836 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1837 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1838 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1839 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1840 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1841 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1842 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1843 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1844 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1845 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1846 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1847 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1848 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1850 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1851 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1852 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1853 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1854 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1855 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1856 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1857 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1858 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1859 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1860 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1861 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1862 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1863 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1864 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1865 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1866 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1867 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1868 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1869 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1870 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1871 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1872 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1873 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764), .A(N14089), .B(N14087), .CI(N14091));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1874 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952), .B(N13727), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1875 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890), .A(N13455), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1876 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1877 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1878 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1879 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1880 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071), .A(N14318), .B(N14316), .CI(N14320));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1881 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146), .B(N14006), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1882 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1883 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1884 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1885 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1886 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1887 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1888 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1889 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1890 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259), .A(N14286), .B(N14284), .CI(N14288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1891 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234), .A(N14160), .B(N14158), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1892 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107), .B(N13849), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_5_I1893 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1894 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1895 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1896 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_5_I1897 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1898 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_5_I1899 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7561));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1900 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I1901 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757), .A(N13455), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1902 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1903 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1904 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1905 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1906 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1907 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1908 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1909 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1910 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1911 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1912 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1913 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1914 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I1918 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1919 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1920 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1921 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046), .A(N14232), .B(N14230), .CI(N14234));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1922 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14]), .A(N13907), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1923 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487), .A(N13735), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15]));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_5_I1924 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1925 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1926 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1927 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1928 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1929 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1930 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390), .A(N14398), .B(N14402), .CI(N14400));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1931 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1932 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1933 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1934 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1935 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125), .B(N14174), .CI(N14178));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1936 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1937 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1938 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15]));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_5_I1939 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1940 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1943 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1944 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1945 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1946 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1947 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1948 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1949 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1950 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1951 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1952 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1953 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1954 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1955 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1956 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13]), .A(N14040), .B(N14038), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1957 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1958 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1959 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1960 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1961 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1962 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1963 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1964 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199), .A(N14326), .B(N14324), .CI(N14328));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1965 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1966 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1967 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14]));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_5_I1968 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1969 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1970 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1971 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1972 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1973 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1974 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1975 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1979 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1980 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1982 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1983 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1984 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1985 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1986 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1987 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]), .A(N14184), .B(N14182), .CI(N14186));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1989 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1990 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1991 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1992 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1993 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329), .A(N14421), .B(N14419), .CI(N14423));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1994 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064), .B(N14278), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1995 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1996 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I1997 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1998 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I1999 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2000 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2001 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2002 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2003 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2004 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2005 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2006 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]), .A(N14294), .B(N14292), .CI(N14296));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2007 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2008 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2009 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2010 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2011 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140), .A(N14384), .B(N14382), .CI(N14386));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2012 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2013 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2014 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2015 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2016 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2017 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2018 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2019 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2020 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2021 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2022 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2023 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2024 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2025 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2026 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]), .A(N14392), .B(N14390), .CI(N14394));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2027 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2028 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2029 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2030 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2031 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2032 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2033 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2034 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2035 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2036 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]), .A(N14471), .B(N14469), .CI(N14473));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2037 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2039 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2040 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2043 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2044 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2045 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2046 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]), .A(N14376), .B(N14374), .CI(N14378));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2047 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2048 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329), .B(N14260), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2049 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2050 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2051 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2052 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2054 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2055 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2056 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2057 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2058 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2059 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2060 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]), .A(N14507), .B(N14505), .CI(N14509));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2061 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2062 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2063 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2066 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2067 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2068 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2069 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2070 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2071 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9]), .CI(N14370));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2072 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2073 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2077 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2078 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2079 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2080 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960), .A(N14456), .B(N14454), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2081 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2082 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2085 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2086 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2087 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2088 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2089 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437), .A(N14489), .B(N14487), .CI(N14491));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2090 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857), .B(N14339), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2091 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2092 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2095 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2096 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2097 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2098 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2099 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592), .A(N14443), .B(N14441), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2104 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2109 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2110 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2111 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2113 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2114 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802), .A(N14481), .B(N14479), .CI(N14483));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2117 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2118 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016), .A(N14517), .B(N14515), .CI(N14519));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2120 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444), .A(N14494), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2122 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2125 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I2130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I2131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936), .A(N14494), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I2133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444), .A1(N14465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I2134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I2136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I2137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I2139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I2140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_5_I2142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_5_I2143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2145 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_5_I2146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I7940 (.Y(N14535), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I7941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558), .A(N14535));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I7942 (.Y(N14543), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I7943 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747), .A(N14543));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I7944 (.Y(N14551), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I7945 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590), .A(N14551));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7807), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7807));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7521), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7521));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7840), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7840));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2161 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2162 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7586), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7586));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7914), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7914));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2166 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7614), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2167 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7614));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2168 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2169 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2170 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7646), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7646));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2172 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2173 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543));
OAI2BB1XL float_div_cynw_cm_float_rcp_E8_M23_5_I2181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749), .A(N12365), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8667 (.Y(N16185), .A(N15293), .B(N12259));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831), .A0N(N15293), .A1N(N12259), .B0(N13254));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8669 (.Y(N16186), .A(N12254));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8670 (.Y(N16199), .A0(N13254), .A1(N16185), .B0(N16186));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8671 (.Y(N16197), .A(N12349));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8672 (.Y(N16203), .A(N16197), .B(N16199));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588), .A0N(N12254), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831), .B0(N12349));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8674 (.Y(N16201), .A(N12249));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8675 (.Y(N16190), .A(N16201), .B(N16203));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8676 (.Y(N16194), .A(N12333));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8677 (.Y(N16193), .A(N16194), .B(N16190));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608), .A(N16193));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899), .A0N(N12244), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608), .B0(N12317));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8657 (.Y(N16169), .A(N12234));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_5_I8658 (.Y(N16171), .AN(N12239), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8659 (.Y(N16168), .A(N16169), .B(N16171));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I8660 (.Y(N16165), .A(N12291), .B(N16168));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8661 (.Y(N16167), .A(N12229));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8662 (.Y(N16173), .A(N16167), .B(N16165));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_5_I8663 (.Y(N16162), .A(N12229), .B(N12291), .C(N16168));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I8664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834), .A(N16171));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I8665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[39]), .A(N16162), .B(N16173));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896), .B(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904));
AO22XL float_div_cynw_cm_float_rcp_E8_M23_5_I2199 (.Y(x[22]), .A0(N12170), .A1(N12164), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[39]), .B1(N12168));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I7938 (.Y(N14526), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834), .B(N12234));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I7939 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38]), .A(N14526));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2201 (.Y(x[21]), .A(N12170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38]), .S0(N12168));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899), .B(N12239));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2203 (.Y(x[20]), .A(N12170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37]), .S0(N12168));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608), .B(N12244));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2205 (.Y(x[19]), .A(N12170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36]), .S0(N12168));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588), .B(N12249));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2207 (.Y(x[18]), .A(N12170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35]), .S0(N12168));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831), .B(N12254));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2209 (.Y(x[17]), .A(N12170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34]), .S0(N12168));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33]), .A(N15293), .B(N12259));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2211 (.Y(x[16]), .A(N12170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33]), .S0(N12168));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32]), .A(N13261), .B(N13263));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2213 (.Y(x[15]), .A(N12170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32]), .S0(N12168));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2215 (.Y(x[14]), .A(N12170), .B(N12266), .S0(N12168));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I7946 (.Y(N14556), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I7947 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30]), .A(N14556));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2217 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[13]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[12]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2221 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[11]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[10]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[9]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[8]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[7]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[6]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[5]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[4]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[3]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[2]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19]), .S0(N11888));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_5_I2240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[1]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18]), .S0(N11888));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I7948 (.Y(N14562), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017));
INVXL float_div_cynw_cm_float_rcp_E8_M23_5_I7949 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17]), .A(N14562));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[0]), .A(N11890), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17]), .S0(N11888));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_5_I2245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_5_I2253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_5_I2254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31]), .AN(a_sign), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29));
EDFFHQX1 x_reg_L0_23__I2278 (.Q(N5677), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_24__I2279 (.Q(N5682), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_25__I2280 (.Q(N5687), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_26__I2281 (.Q(N5692), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_27__I2282 (.Q(N5697), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_28__I2283 (.Q(N5702), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_29__I2284 (.Q(N5707), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_30__I2285 (.Q(N5712), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_31__I2286 (.Q(N5717), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_0__I2287 (.Q(x[0]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_1__I2288 (.Q(x[1]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_2__I2289 (.Q(x[2]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_3__I2290 (.Q(x[3]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_4__I2291 (.Q(x[4]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_5__I2292 (.Q(x[5]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_6__I2293 (.Q(x[6]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_7__I2294 (.Q(x[7]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_8__I2295 (.Q(x[8]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_9__I2296 (.Q(x[9]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__I2297 (.Q(x[10]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_11__I2298 (.Q(x[11]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__I2299 (.Q(x[12]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__I2310 (.Q(x[23]), .D(N5677), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_24__I2311 (.Q(x[24]), .D(N5682), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_25__I2312 (.Q(x[25]), .D(N5687), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_26__I2313 (.Q(x[26]), .D(N5692), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_27__I2314 (.Q(x[27]), .D(N5697), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_28__I2315 (.Q(x[28]), .D(N5702), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_29__I2316 (.Q(x[29]), .D(N5707), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_30__I2317 (.Q(x[30]), .D(N5712), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_31__I2318 (.Q(x[31]), .D(N5717), .E(bdw_enable), .CK(aclk));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[14] = x[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[15] = x[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[19] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[20] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[16] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  srD0Tgzcqhw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



