/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:40:44 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_2_1 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__9,
	inst_cellmath__10,
	inst_cellmath__11,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__16,
	inst_cellmath__17,
	inst_cellmath__18;
wire [8:0] inst_cellmath__27;
wire [7:0] inst_cellmath__29;
wire  inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__32;
wire [49:0] inst_cellmath__33;
wire [7:0] inst_cellmath__35;
wire [49:0] inst_cellmath__36,
	inst_cellmath__37;
wire [25:0] inst_cellmath__39;
wire  inst_cellmath__42,
	inst_cellmath__43,
	inst_cellmath__44;
wire [26:0] inst_cellmath__45;
wire  inst_cellmath__48;
wire [5:0] inst_cellmath__49;
wire [24:0] inst_cellmath__50;
wire  inst_cellmath__53,
	inst_cellmath__54,
	inst_cellmath__55;
wire [23:0] inst_cellmath__57;
wire [9:0] inst_cellmath__59;
wire  inst_cellmath__62,
	inst_cellmath__63;
wire [22:0] inst_cellmath__64;
wire  inst_cellmath__66;
wire [7:0] inst_cellmath__68;
wire  inst_cellmath__70,
	inst_cellmath__71;
wire N547,N556,N557,N558,N559,N560,N561 
	,N562,N563,N566,N568,N569,N570,N571,N572 
	,N574,N575,N626,N627,N628,N630,N634,N635 
	,N636,N639,N645,N650,N651,N652,N653,N655 
	,N656,N657,N658,N659,N660,N661,N662,N663 
	,N664,N665,N666,N667,N668,N669,N670,N671 
	,N672,N673,N674,N675,N676,N677,N706,N710 
	,N3083,N3085,N3106,N3114,N3117,N3119,N3123,N3125 
	,N3128,N3134,N3138,N3168,N3170,N3191,N3199,N3202 
	,N3204,N3208,N3210,N3213,N3219,N3223,N3319,N3321 
	,N3327,N3330,N3331,N3333,N3337,N3338,N3343,N3348 
	,N3358,N3362,N3364,N3367,N3459,N3494,N3597,N3604 
	,N3612,N3614,N3617,N3620,N3627,N3655,N3656,N3695 
	,N3766,N3768,N3769,N3770,N3772,N3774,N3775,N3777 
	,N3778,N3779,N3781,N3783,N3784,N3785,N3786,N3788 
	,N3790,N3792,N3793,N3794,N3795,N3798,N3800,N3802 
	,N3803,N3805,N3807,N3809,N3810,N3811,N3812,N3815 
	,N3816,N3817,N3819,N3821,N3822,N3823,N3825,N3827 
	,N3828,N3830,N3832,N3833,N3835,N3837,N3839,N3840 
	,N3841,N3842,N3845,N3846,N3847,N3849,N3851,N3852 
	,N3853,N3854,N3856,N3858,N3860,N3861,N3863,N3865 
	,N3866,N3868,N3871,N3873,N3875,N3876,N3877,N3878 
	,N3880,N3882,N3884,N3885,N3886,N3888,N3890,N3891 
	,N3892,N3894,N3896,N3897,N3899,N3901,N3903,N3904 
	,N3905,N3906,N3909,N3910,N3911,N3912,N3914,N3916 
	,N3918,N3919,N3920,N3922,N3924,N3925,N3927,N3929 
	,N3931,N3932,N3933,N3934,N3937,N3938,N3940,N3942 
	,N3943,N3944,N3945,N3947,N3948,N3950,N3952,N3953 
	,N3955,N3957,N3958,N3959,N3960,N3961,N3963,N3966 
	,N3967,N3968,N3970,N3972,N3973,N3974,N3975,N3977 
	,N3979,N3982,N3983,N4205,N4261,N4265,N4271,N4274 
	,N4279,N4282,N4291,N4294,N4300,N4328,N4508,N4510 
	,N4511,N4512,N4518,N4521,N4524,N4529,N4530,N4533 
	,N4534,N4537,N4539,N4540,N4541,N4544,N4546,N4549 
	,N4550,N4554,N4556,N4558,N4561,N4562,N4564,N4566 
	,N4568,N4572,N4575,N4576,N4581,N4582,N4585,N4586 
	,N4588,N4589,N4592,N4593,N4594,N4599,N4601,N4604 
	,N4605,N4609,N4614,N4617,N4618,N4622,N4623,N4629 
	,N4630,N4631,N4712,N4714,N4715,N4716,N4717,N4719 
	,N4720,N4723,N4724,N4725,N4726,N4728,N4729,N4730 
	,N4733,N4734,N4735,N4736,N4738,N4740,N4743,N4744 
	,N4745,N4747,N4748,N4750,N4751,N4752,N4754,N4756 
	,N4757,N4758,N4760,N4761,N4762,N4765,N4766,N4768 
	,N4769,N4771,N4773,N4775,N4776,N4777,N4779,N4780 
	,N4781,N4782,N4784,N4786,N4788,N4789,N4790,N4792 
	,N4793,N4795,N4797,N4798,N4799,N4801,N4802,N4805 
	,N4806,N4931,N4952,N5001,N5004,N5010,N5016,N5017 
	,N5019,N5020,N5022,N5023,N5025,N5026,N5029,N5030 
	,N5031,N5033,N5034,N5036,N5037,N5038,N5040,N5042 
	,N5043,N5045,N5047,N5049,N5050,N5052,N5053,N5054 
	,N5056,N5057,N5059,N5060,N5062,N5063,N5065,N5066 
	,N5068,N5069,N5071,N5072,N5074,N5076,N5077,N5079 
	,N5080,N5081,N5083,N5084,N5086,N5087,N5090,N5092 
	,N5093,N5094,N5096,N5098,N5099,N5101,N5102,N5104 
	,N5105,N5106,N5108,N5109,N5111,N5113,N5114,N5116 
	,N5117,N5119,N5121,N5123,N5124,N5126,N5127,N5128 
	,N5130,N5131,N5133,N5135,N5136,N5138,N5139,N5141 
	,N5142,N5143,N5145,N5146,N5148,N5149,N5151,N5153 
	,N5154,N5155,N5157,N5158,N5160,N5162,N5163,N5164 
	,N5166,N5167,N5169,N5171,N5172,N5173,N5175,N5176 
	,N5178,N5179,N5354,N5374,N5418,N5421,N5426,N5428 
	,N5429,N5434,N5436,N5438,N5445,N5446,N5449,N5452 
	,N5454,N5456,N5461,N5464,N5466,N5473,N5474,N5477 
	,N5480,N5482,N5580,N5583,N5584,N5592,N5600,N5605 
	,N5610,N5612,N5614,N5617,N5619,N5622,N5630,N5733 
	,N5745,N5751,N5769,N5790,N5796,N5801,N5804,N5808 
	,N5812,N5817,N5820,N5821,N5825,N5831,N5834,N5839 
	,N5844,N5847,N5851,N5856,N5860,N5864,N5868,N5873 
	,N5875,N5877,N5881,N5886,N5889,N7112,N7129,N7134 
	,N7135,N7138,N7139,N7140,N7141,N7143,N7149,N7157 
	,N11648,N11649,N11650,N11651,N11652,N11653,N11788,N11789 
	,N11950,N11972,N11973,N11975,N11977,N11980,N11981,N11985 
	,N11986,N12004,N12005,N12016,N12017,N12033,N12036,N12038 
	,N12040,N12043,N12046,N12049,N12052,N12054,N12057,N12060 
	,N12062,N12063,N12066,N12070,N12073,N12075,N12076,N12079 
	,N12083,N12086,N12088,N12091,N12092,N12123,N12125,N12129 
	,N12134,N12139,N12145,N12148,N12151,N12157,N12160,N12162 
	,N12165,N12174,N12177,N12184,N12188,N12189,N12194,N12241 
	,N12252,N12264,N12275,N12287,N12298,N12310,N12314,N12317 
	,N12319,N12321,N12323,N12333,N12336,N12338,N12339,N12341 
	,N12343,N12344,N12346,N12347,N12350,N12351,N12352,N12368 
	,N12369,N12371,N12373,N12374,N12375,N12378,N12379,N12380 
	,N12382,N12384,N12386,N12387,N12389,N12391,N12409,N12410 
	,N12412,N12414,N12415,N12416,N12419,N12420,N12421,N12423 
	,N12425,N12427,N12428,N12430,N12432,N12450,N12451,N12453 
	,N12455,N12456,N12457,N12460,N12461,N12462,N12464,N12466 
	,N12468,N12469,N12471,N12473,N12492,N12499,N12507,N12518 
	,N12547,N12548,N12550,N12557,N12558,N12560,N12565,N12567 
	,N12573,N12575,N12578,N12582,N12585,N12592,N12595,N12633 
	,N12635,N12638,N12639,N12642,N12650,N12652,N12658,N12661 
	,N12662,N12687,N12695,N12699,N12706,N12713,N12720,N12727 
	,N12734,N12741,N12748,N12755;
XOR2XL cynw_cm_float_add2_ieee_I462 (.Y(inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
NAND2XL inst_cellmath__9_0_I463 (.Y(N3083), .A(a_exp[0]), .B(a_exp[1]));
AND4XL inst_cellmath__9_0_I7167 (.Y(N3085), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I2721 (.Y(N7149), .A(a_exp[7]), .B(a_exp[6]), .C(N3085));
NOR2XL hyperpropagate_4_1_A_I2722 (.Y(inst_cellmath__9), .A(N3083), .B(N7149));
NOR2XL inst_cellmath__10__1__I476 (.Y(N3106), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__10__1__I477 (.Y(N3114), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__10__1__I478 (.Y(N3125), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__10__1__I479 (.Y(N3134), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__10__1__I7168 (.Y(N3119), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__10__1__I7169 (.Y(N3128), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__10__1__I7170 (.Y(N3138), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
INVXL inst_cellmath__64__48__2WWMM_I6635 (.Y(N11652), .A(a_man[0]));
INVXL cynw_cm_float_add2_ieee_I7099 (.Y(N11653), .A(N11652));
NOR4X1 inst_cellmath__10__1__I483 (.Y(N3123), .A(N11653), .B(a_man[1]), .C(a_man[2]), .D(N3119));
NAND4XL inst_cellmath__10__1__I485 (.Y(N3117), .A(N3106), .B(N3125), .C(N3114), .D(N3134));
NOR4BX1 inst_cellmath__10__1__I7171 (.Y(inst_cellmath__10), .AN(N3123), .B(N3117), .C(N3128), .D(N3138));
NAND2XL inst_cellmath__14_0_I489 (.Y(N3168), .A(b_exp[0]), .B(b_exp[1]));
AND4XL inst_cellmath__14_0_I7172 (.Y(N3170), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL hyperpropagate_4_1_A_I2723 (.Y(N7157), .A(b_exp[7]), .B(b_exp[6]), .C(N3170));
NOR2XL hyperpropagate_4_1_A_I2724 (.Y(inst_cellmath__14), .A(N3168), .B(N7157));
NOR2XL inst_cellmath__15__3__I502 (.Y(N3191), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__15__3__I503 (.Y(N3199), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__15__3__I504 (.Y(N3210), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__15__3__I505 (.Y(N3219), .A(b_man[4]), .B(b_man[3]));
OR4X1 inst_cellmath__15__3__I7173 (.Y(N3204), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__15__3__I7174 (.Y(N3213), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__15__3__I7175 (.Y(N3223), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4X1 inst_cellmath__15__3__I509 (.Y(N3208), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N3204));
NAND4XL inst_cellmath__15__3__I511 (.Y(N3202), .A(N3191), .B(N3210), .C(N3199), .D(N3219));
NOR4BX1 inst_cellmath__15__3__I7176 (.Y(inst_cellmath__15), .AN(N3208), .B(N3202), .C(N3213), .D(N3223));
AND2XL inst_cellmath__62_0_I6929 (.Y(inst_cellmath__17), .A(inst_cellmath__14), .B(inst_cellmath__15));
AND2XL inst_cellmath__62_0_I6928 (.Y(inst_cellmath__12), .A(inst_cellmath__9), .B(inst_cellmath__10));
AND3XL cynw_cm_float_add2_ieee_I515 (.Y(N547), .A(inst_cellmath__17), .B(inst_cellmath__12), .C(inst_cellmath__39[25]));
NOR2BX1 cynw_cm_float_add2_ieee_I516 (.Y(inst_cellmath__13), .AN(inst_cellmath__9), .B(inst_cellmath__10));
NOR2BX1 cynw_cm_float_add2_ieee_I517 (.Y(inst_cellmath__18), .AN(inst_cellmath__14), .B(inst_cellmath__15));
OR4X1 cynw_cm_float_add2_ieee_I7177 (.Y(N12062), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 cynw_cm_float_add2_ieee_I7178 (.Y(N12075), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL cynw_cm_float_add2_ieee_I6901 (.Y(inst_cellmath__11), .A(N12062), .B(N12075));
OR4X1 cynw_cm_float_add2_ieee_I7179 (.Y(N12040), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 cynw_cm_float_add2_ieee_I7180 (.Y(N12054), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL cynw_cm_float_add2_ieee_I6904 (.Y(inst_cellmath__16), .A(N12040), .B(N12054));
INVX1 cynw_cm_float_add2_ieee_I15 (.Y(N556), .A(b_exp[0]));
INVXL cynw_cm_float_add2_ieee_I16 (.Y(N557), .A(b_exp[1]));
INVXL cynw_cm_float_add2_ieee_I17 (.Y(N558), .A(b_exp[2]));
INVXL cynw_cm_float_add2_ieee_I18 (.Y(N559), .A(b_exp[3]));
INVXL cynw_cm_float_add2_ieee_I19 (.Y(N560), .A(b_exp[4]));
INVXL cynw_cm_float_add2_ieee_I20 (.Y(N561), .A(b_exp[5]));
ADDHX1 cynw_cm_float_add2_ieee_I6886 (.CO(N3321), .S(N12017), .A(N556), .B(a_exp[0]));
ADDFX1 inst_cellmath__28__8__I536 (.CO(N3364), .S(N566), .A(N557), .B(a_exp[1]), .CI(N3321));
ADDFX1 cynw_cm_float_add2_ieee_I7094 (.CO(N3338), .S(N12518), .A(a_exp[2]), .B(N3364), .CI(N558));
ADDFX1 inst_cellmath__28__8__I538 (.CO(N3358), .S(N568), .A(N559), .B(a_exp[3]), .CI(N3338));
ADDFX1 inst_cellmath__28__8__I539 (.CO(N3331), .S(N569), .A(N560), .B(a_exp[4]), .CI(N3358));
OR2XL inst_cellmath__28__8__I545 (.Y(N3333), .A(a_exp[0]), .B(N556));
ADDFX1 inst_cellmath__28__8__I546 (.CO(N3327), .S(inst_cellmath__27[1]), .A(N557), .B(a_exp[1]), .CI(N3333));
ADDFX1 inst_cellmath__28__8__I547 (.CO(N3348), .S(inst_cellmath__27[2]), .A(N558), .B(a_exp[2]), .CI(N3327));
ADDFX1 inst_cellmath__28__8__I548 (.CO(N3319), .S(inst_cellmath__27[3]), .A(N559), .B(a_exp[3]), .CI(N3348));
ADDFX1 inst_cellmath__28__8__I549 (.CO(N3343), .S(inst_cellmath__27[4]), .A(N560), .B(a_exp[4]), .CI(N3319));
ADDFX1 inst_cellmath__28__8__I550 (.CO(N3362), .S(inst_cellmath__27[5]), .A(N561), .B(a_exp[5]), .CI(N3343));
INVXL inst_cellmath__34_0_I7150 (.Y(N562), .A(b_exp[6]));
ADDFX1 inst_cellmath__28__8__I551 (.CO(N3337), .S(inst_cellmath__27[6]), .A(N562), .B(a_exp[6]), .CI(N3362));
INVXL inst_cellmath__34_0_I7151 (.Y(N563), .A(b_exp[7]));
ADDFX1 inst_cellmath__28__8__I552 (.CO(N3330), .S(inst_cellmath__27[7]), .A(N563), .B(a_exp[7]), .CI(N3337));
INVX2 inst_cellmath__34_0_I563 (.Y(N3459), .A(a_man[20]));
INVX2 inst_cellmath__34_0_I6874 (.Y(N11986), .A(a_man[2]));
CLKINVX6 inst_cellmath__34_0_I6875 (.Y(N11981), .A(b_man[0]));
NOR2X6 inst_cellmath__34_0_I6876 (.Y(N11977), .A(a_man[0]), .B(N11981));
INVX8 inst_cellmath__34_0_I6877 (.Y(N11980), .A(a_man[1]));
NOR2X4 inst_cellmath__34_0_I6878 (.Y(N11985), .A(b_man[1]), .B(N11980));
AOI21X4 inst_cellmath__34_0_I6879 (.Y(N11972), .A0(b_man[1]), .A1(N11980), .B0(N11977));
INVX1 inst_cellmath__34_0_I6880 (.Y(N11975), .A(b_man[2]));
NOR2X4 inst_cellmath__34_0_I6882 (.Y(N11973), .A(b_man[2]), .B(N11986));
INVX2 inst_cellmath__34_0_I6986 (.Y(N12319), .A(a_man[6]));
INVX2 inst_cellmath__34_0_I6987 (.Y(N12323), .A(b_man[5]));
INVX2 inst_cellmath__34_0_I6988 (.Y(N12310), .A(b_man[7]));
INVXL inst_cellmath__34_0_I7029 (.Y(N12346), .A(a_man[4]));
INVXL inst_cellmath__34_0_I7030 (.Y(N12351), .A(b_man[3]));
INVX2 inst_cellmath__34_0_I7031 (.Y(N12344), .A(a_man[3]));
NOR2BX1 inst_cellmath__34_0_I7032 (.Y(N12347), .AN(N12351), .B(N12344));
NOR2BX2 inst_cellmath__34_0_I7033 (.Y(N12338), .AN(N12344), .B(N12351));
NOR2X2 inst_cellmath__34_0_I7034 (.Y(N12339), .A(N11975), .B(a_man[2]));
NOR3X6 inst_cellmath__34_0_I7035 (.Y(N12343), .A(N11985), .B(N11973), .C(N11972));
NOR3X4 inst_cellmath__34_0_I7036 (.Y(N12352), .A(N12339), .B(N12338), .C(N12343));
INVXL inst_cellmath__34_0_I7037 (.Y(N12333), .A(b_man[4]));
NOR2BX1 inst_cellmath__34_0_I7038 (.Y(N12336), .AN(N12346), .B(N12333));
NOR2BX1 inst_cellmath__34_0_I7039 (.Y(N12350), .AN(N12333), .B(N12346));
NOR3X2 inst_cellmath__34_0_I7040 (.Y(N12341), .A(N12347), .B(N12350), .C(N12352));
NOR2X2 inst_cellmath__34_0_I7041 (.Y(N12314), .A(N12336), .B(N12341));
ACHCONX2 inst_cellmath__34_0_I6990 (.CON(N12317), .A(N12323), .B(a_man[5]), .CI(N12314));
ACHCONX2 inst_cellmath__34_0_I6991 (.CON(N12321), .A(N12319), .B(b_man[6]), .CI(N12317));
INVXL inst_cellmath__34_0_I7077 (.Y(N12468), .A(a_man[10]));
INVXL inst_cellmath__34_0_I7078 (.Y(N12451), .A(b_man[9]));
INVXL inst_cellmath__34_0_I7079 (.Y(N12461), .A(b_man[8]));
NAND2X1 inst_cellmath__34_0_I7080 (.Y(N12456), .A(N12461), .B(a_man[8]));
INVX1 inst_cellmath__34_0_I7081 (.Y(N12453), .A(a_man[9]));
NOR2BX1 inst_cellmath__34_0_I7082 (.Y(N12457), .AN(N12451), .B(N12453));
INVXL inst_cellmath__34_0_I7083 (.Y(N12450), .A(N12451));
INVXL inst_cellmath__34_0_I7084 (.Y(N12460), .A(N12461));
INVX1 inst_cellmath__34_0_I7085 (.Y(N12466), .A(a_man[8]));
ACHCONX2 inst_cellmath__34_0_I7086 (.CON(N12471), .A(N12310), .B(a_man[7]), .CI(N12321));
AOI222X4 inst_cellmath__34_0_I7087 (.Y(N12462), .A0(N12460), .A1(N12466), .B0(N12453), .B1(N12450), .C0(N12456), .C1(N12471));
INVXL inst_cellmath__34_0_I7088 (.Y(N12469), .A(b_man[10]));
NOR2BX1 inst_cellmath__34_0_I7089 (.Y(N12473), .AN(N12468), .B(N12469));
NOR2BX1 inst_cellmath__34_0_I7090 (.Y(N12464), .AN(N12469), .B(N12468));
NOR3X4 inst_cellmath__34_0_I7091 (.Y(N12455), .A(N12464), .B(N12457), .C(N12462));
NOR2X4 inst_cellmath__34_0_I7092 (.Y(N12298), .A(N12473), .B(N12455));
INVX2 inst_cellmath__34_0_I6980 (.Y(N12287), .A(b_man[11]));
INVXL inst_cellmath__34_0_I7060 (.Y(N12427), .A(a_man[14]));
INVXL inst_cellmath__34_0_I7061 (.Y(N12410), .A(b_man[13]));
INVXL inst_cellmath__34_0_I7062 (.Y(N12419), .A(b_man[12]));
NAND2XL inst_cellmath__34_0_I7063 (.Y(N12415), .A(N12419), .B(a_man[12]));
INVXL inst_cellmath__34_0_I7064 (.Y(N12412), .A(a_man[13]));
NOR2BX1 inst_cellmath__34_0_I7065 (.Y(N12416), .AN(N12410), .B(N12412));
INVXL inst_cellmath__34_0_I7066 (.Y(N12409), .A(N12410));
INVXL inst_cellmath__34_0_I7067 (.Y(N12420), .A(N12419));
INVXL inst_cellmath__34_0_I7068 (.Y(N12425), .A(a_man[12]));
ACHCONX2 inst_cellmath__34_0_I7069 (.CON(N12430), .A(a_man[11]), .B(N12287), .CI(N12298));
AOI222X4 inst_cellmath__34_0_I7070 (.Y(N12421), .A0(N12420), .A1(N12425), .B0(N12412), .B1(N12409), .C0(N12415), .C1(N12430));
INVXL inst_cellmath__34_0_I7071 (.Y(N12428), .A(b_man[14]));
NOR2BX1 inst_cellmath__34_0_I7072 (.Y(N12432), .AN(N12427), .B(N12428));
NOR2BX1 inst_cellmath__34_0_I7073 (.Y(N12423), .AN(N12428), .B(N12427));
NOR3X4 inst_cellmath__34_0_I7074 (.Y(N12414), .A(N12423), .B(N12416), .C(N12421));
NOR2X4 inst_cellmath__34_0_I7075 (.Y(N12275), .A(N12432), .B(N12414));
INVX2 inst_cellmath__34_0_I6972 (.Y(N12264), .A(b_man[15]));
INVXL inst_cellmath__34_0_I7043 (.Y(N12386), .A(a_man[18]));
INVXL inst_cellmath__34_0_I7044 (.Y(N12369), .A(b_man[17]));
INVXL inst_cellmath__34_0_I7045 (.Y(N12378), .A(b_man[16]));
NAND2XL inst_cellmath__34_0_I7046 (.Y(N12374), .A(N12378), .B(a_man[16]));
INVXL inst_cellmath__34_0_I7047 (.Y(N12371), .A(a_man[17]));
NOR2BX1 inst_cellmath__34_0_I7048 (.Y(N12375), .AN(N12369), .B(N12371));
INVXL inst_cellmath__34_0_I7049 (.Y(N12368), .A(N12369));
INVXL inst_cellmath__34_0_I7050 (.Y(N12379), .A(N12378));
INVX1 inst_cellmath__34_0_I7051 (.Y(N12384), .A(a_man[16]));
ACHCONX2 inst_cellmath__34_0_I7052 (.CON(N12389), .A(N12264), .B(a_man[15]), .CI(N12275));
AOI222X4 inst_cellmath__34_0_I7053 (.Y(N12380), .A0(N12379), .A1(N12384), .B0(N12371), .B1(N12368), .C0(N12374), .C1(N12389));
INVXL inst_cellmath__34_0_I7054 (.Y(N12387), .A(b_man[18]));
NOR2BX1 inst_cellmath__34_0_I7055 (.Y(N12391), .AN(N12386), .B(N12387));
NOR2BX1 inst_cellmath__34_0_I7056 (.Y(N12382), .AN(N12387), .B(N12386));
NOR3X4 inst_cellmath__34_0_I7057 (.Y(N12373), .A(N12382), .B(N12375), .C(N12380));
NOR2X4 inst_cellmath__34_0_I7058 (.Y(N12252), .A(N12391), .B(N12373));
INVX2 inst_cellmath__34_0_I6964 (.Y(N12241), .A(b_man[19]));
ACHCONX2 inst_cellmath__34_0_I6968 (.CON(N3494), .A(N12241), .B(a_man[19]), .CI(N12252));
INVXL inst_cellmath__34_0_I7156 (.Y(N11950), .A(b_man[21]));
ADDFX1 inst_cellmath__34_0_I7152 (.CO(N12635), .S(N570), .A(a_exp[5]), .B(N561), .CI(N3331));
ADDFX1 inst_cellmath__34_0_I7153 (.CO(N12652), .S(N571), .A(a_exp[6]), .B(N562), .CI(N12635));
ADDFX1 inst_cellmath__34_0_I7154 (.CO(N3367), .S(N572), .A(N563), .B(a_exp[7]), .CI(N12652));
INVXL inst_cellmath__34_0_I7155 (.Y(N12638), .A(a_man[22]));
AND2XL inst_cellmath__34_0_I7185 (.Y(N12662), .A(N12638), .B(b_man[22]));
NAND2XL inst_cellmath__34_0_I7160 (.Y(N12633), .A(a_man[21]), .B(N11950));
OR2XL inst_cellmath__34_0_I7186 (.Y(N12642), .A(a_man[21]), .B(N11950));
ACHCONX2 inst_cellmath__34_0_I7162 (.CON(N12650), .A(N3459), .B(b_man[20]), .CI(N3494));
NAND2X4 inst_cellmath__34_0_I7163 (.Y(N12658), .A(N12642), .B(N12650));
OR2XL inst_cellmath__34_0_I7188 (.Y(N12661), .A(b_man[22]), .B(N12638));
AOI31X4 inst_cellmath__34_0_I7165 (.Y(N12639), .A0(N12661), .A1(N12633), .A2(N12658), .B0(N12662));
NOR2X4 inst_cellmath__34_0_I7166 (.Y(N575), .A(N3367), .B(N12639));
CLKINVX8 cynw_cm_float_add2_ieee_I7096 (.Y(inst_cellmath__27[8]), .A(N3330));
INVXL inst_cellmath__35_0_I625 (.Y(N3617), .A(inst_cellmath__27[1]));
INVXL inst_cellmath__35_0_I627 (.Y(N3597), .A(inst_cellmath__27[3]));
INVXL inst_cellmath__35_0_I628 (.Y(N3604), .A(inst_cellmath__27[4]));
INVXL inst_cellmath__35_0_I629 (.Y(N3612), .A(inst_cellmath__27[5]));
INVXL inst_cellmath__35_0_I630 (.Y(N3620), .A(inst_cellmath__27[6]));
INVXL inst_cellmath__35_0_I631 (.Y(N3627), .A(inst_cellmath__27[7]));
INVX1 cynw_cm_float_add2_ieee_I7097 (.Y(N3614), .A(inst_cellmath__27[8]));
AOI22X1 inst_cellmath__35_0_I634 (.Y(inst_cellmath__35[1]), .A0(N3617), .A1(N3614), .B0(N566), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I636 (.Y(inst_cellmath__35[3]), .A0(N3614), .A1(N3597), .B0(N568), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I637 (.Y(inst_cellmath__35[4]), .A0(N3614), .A1(N3604), .B0(N569), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I638 (.Y(inst_cellmath__35[5]), .A0(N3614), .A1(N3612), .B0(N570), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I639 (.Y(inst_cellmath__35[6]), .A0(N3614), .A1(N3620), .B0(N571), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I640 (.Y(inst_cellmath__35[7]), .A0(N3614), .A1(N3627), .B0(N572), .B1(inst_cellmath__27[8]));
INVXL cynw_cm_float_add2_ieee_I7095 (.Y(N12499), .A(inst_cellmath__27[2]));
AOI22XL cynw_cm_float_add2_ieee_I7098 (.Y(inst_cellmath__35[2]), .A0(N12518), .A1(inst_cellmath__27[8]), .B0(N12499), .B1(N3614));
OAI211X1 inst_cellmath__30_0_I641 (.Y(N3656), .A0(inst_cellmath__35[2]), .A1(inst_cellmath__35[1]), .B0(inst_cellmath__35[4]), .C0(inst_cellmath__35[3]));
NOR3BXL inst_cellmath__30_0_I642 (.Y(N3655), .AN(N3656), .B(inst_cellmath__35[6]), .C(inst_cellmath__35[5]));
NAND2BX1 inst_cellmath__30_0_I643 (.Y(inst_cellmath__30), .AN(inst_cellmath__35[7]), .B(N3655));
NOR2X6 cynw_cm_float_add2_ieee_I7118 (.Y(inst_cellmath__32), .A(inst_cellmath__27[8]), .B(N575));
INVX12 cynw_cm_float_add2_ieee_I7100 (.Y(N3695), .A(inst_cellmath__32));
MX2XL cynw_cm_float_add2_ieee_I649 (.Y(inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I650 (.Y(inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I653 (.Y(inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I654 (.Y(inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I655 (.Y(inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I656 (.Y(inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I657 (.Y(inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I658 (.Y(inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I659 (.Y(inst_cellmath__36[37]), .A(b_man[11]), .B(a_man[11]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I660 (.Y(inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I661 (.Y(inst_cellmath__36[39]), .A(b_man[13]), .B(a_man[13]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I662 (.Y(inst_cellmath__36[40]), .A(b_man[14]), .B(a_man[14]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I663 (.Y(inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I664 (.Y(inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I665 (.Y(inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I666 (.Y(inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(N3695));
XOR2XL cynw_cm_float_add2_ieee_I6887 (.Y(N12005), .A(N556), .B(a_exp[0]));
MX2XL cynw_cm_float_add2_ieee_I7101 (.Y(inst_cellmath__36[26]), .A(b_man[0]), .B(N11653), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I7102 (.Y(inst_cellmath__36[29]), .A(b_man[3]), .B(a_man[3]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I7103 (.Y(inst_cellmath__36[30]), .A(b_man[4]), .B(a_man[4]), .S0(N3695));
AOI22XL cynw_cm_float_add2_ieee_I7104 (.Y(N12492), .A0(N12017), .A1(inst_cellmath__27[8]), .B0(N12005), .B1(N3614));
INVX1 cynw_cm_float_add2_ieee_I7105 (.Y(N3947), .A(N12492));
MX2XL cynw_cm_float_add2_ieee_I7108 (.Y(N3841), .A(inst_cellmath__36[30]), .B(inst_cellmath__36[29]), .S0(N3947));
CLKINVX6 cynw_cm_float_add2_ieee_I7109 (.Y(N3777), .A(inst_cellmath__35[2]));
CLKINVX6 cynw_cm_float_add2_ieee_I7110 (.Y(N3827), .A(N3777));
NAND2XL hyperpropagate_3_1_A_I7319 (.Y(N12687), .A(inst_cellmath__36[26]), .B(N3777));
NOR2XL hyperpropagate_3_1_A_I7320 (.Y(N12507), .A(N3947), .B(N12687));
AOI21X1 cynw_cm_float_add2_ieee_I7113 (.Y(N3909), .A0(N3827), .A1(N3841), .B0(N12507));
MXI2XL cynw_cm_float_add2_ieee_I6893 (.Y(N12004), .A(b_man[20]), .B(a_man[20]), .S0(N3695));
MXI2X1 cynw_cm_float_add2_ieee_I6894 (.Y(N12016), .A(b_man[19]), .B(a_man[19]), .S0(N3695));
MXI2XL cynw_cm_float_add2_ieee_I6895 (.Y(N3943), .A(N12004), .B(N12016), .S0(N3947));
INVXL cynw_cm_float_add2_ieee_I6896 (.Y(inst_cellmath__36[45]), .A(N12016));
INVXL cynw_cm_float_add2_ieee_I6897 (.Y(inst_cellmath__36[46]), .A(N12004));
MX2XL cynw_cm_float_add2_ieee_I669 (.Y(inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(N3695));
MX2XL cynw_cm_float_add2_ieee_I670 (.Y(inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(N3695));
MX2XL inst_cellmath__37_0_I673 (.Y(N3911), .A(inst_cellmath__36[27]), .B(inst_cellmath__36[26]), .S0(N3947));
MX2X1 inst_cellmath__37_0_I674 (.Y(N3959), .A(inst_cellmath__36[28]), .B(inst_cellmath__36[27]), .S0(N3947));
MX2XL inst_cellmath__37_0_I675 (.Y(N3793), .A(inst_cellmath__36[29]), .B(inst_cellmath__36[28]), .S0(N3947));
MX2XL inst_cellmath__37_0_I677 (.Y(N3885), .A(inst_cellmath__36[31]), .B(inst_cellmath__36[30]), .S0(N3947));
MX2XL inst_cellmath__37_0_I678 (.Y(N3932), .A(inst_cellmath__36[32]), .B(inst_cellmath__36[31]), .S0(N3947));
MX2XL inst_cellmath__37_0_I679 (.Y(N3983), .A(inst_cellmath__36[33]), .B(inst_cellmath__36[32]), .S0(N3947));
MX2X1 inst_cellmath__37_0_I680 (.Y(N3810), .A(inst_cellmath__36[34]), .B(inst_cellmath__36[33]), .S0(N3947));
MX2XL inst_cellmath__37_0_I681 (.Y(N3861), .A(inst_cellmath__36[35]), .B(inst_cellmath__36[34]), .S0(N3947));
MX2X1 inst_cellmath__37_0_I682 (.Y(N3905), .A(inst_cellmath__36[36]), .B(inst_cellmath__36[35]), .S0(N3947));
MX2XL inst_cellmath__37_0_I683 (.Y(N3953), .A(inst_cellmath__36[37]), .B(inst_cellmath__36[36]), .S0(N3947));
MX2XL inst_cellmath__37_0_I684 (.Y(N3784), .A(inst_cellmath__36[38]), .B(inst_cellmath__36[37]), .S0(N3947));
MX2XL inst_cellmath__37_0_I685 (.Y(N3833), .A(inst_cellmath__36[39]), .B(inst_cellmath__36[38]), .S0(N3947));
MX2XL inst_cellmath__37_0_I686 (.Y(N3876), .A(inst_cellmath__36[40]), .B(inst_cellmath__36[39]), .S0(N3947));
MX2X1 inst_cellmath__37_0_I687 (.Y(N3925), .A(inst_cellmath__36[41]), .B(inst_cellmath__36[40]), .S0(N3947));
MX2XL inst_cellmath__37_0_I688 (.Y(N3973), .A(inst_cellmath__36[42]), .B(inst_cellmath__36[41]), .S0(N3947));
MX2XL inst_cellmath__37_0_I689 (.Y(N3803), .A(inst_cellmath__36[43]), .B(inst_cellmath__36[42]), .S0(N3947));
MX2XL inst_cellmath__37_0_I690 (.Y(N3852), .A(inst_cellmath__36[44]), .B(inst_cellmath__36[43]), .S0(N3947));
MX2XL inst_cellmath__37_0_I691 (.Y(N3897), .A(inst_cellmath__36[45]), .B(inst_cellmath__36[44]), .S0(N3947));
MX2XL inst_cellmath__37_0_I693 (.Y(N3775), .A(inst_cellmath__36[47]), .B(inst_cellmath__36[46]), .S0(N3947));
MX2XL inst_cellmath__37_0_I694 (.Y(N3822), .A(inst_cellmath__36[48]), .B(inst_cellmath__36[47]), .S0(N3947));
NAND2BXL inst_cellmath__37_0_I695 (.Y(N3868), .AN(inst_cellmath__36[48]), .B(N3947));
NAND3BXL inst_cellmath__37_0_I7192 (.Y(N3966), .AN(N3947), .B(inst_cellmath__36[26]), .C(N3827));
NAND2XL inst_cellmath__37_0_I699 (.Y(N3845), .A(N3827), .B(N3911));
NAND2XL inst_cellmath__37_0_I700 (.Y(N3937), .A(N3827), .B(N3959));
NAND2XL inst_cellmath__37_0_I701 (.Y(N3815), .A(N3827), .B(N3793));
AOI22X1 inst_cellmath__37_0_I703 (.Y(N3957), .A0(N3827), .A1(N3885), .B0(N3911), .B1(N3777));
AOI22X1 inst_cellmath__37_0_I704 (.Y(N3790), .A0(N3827), .A1(N3932), .B0(N3959), .B1(N3777));
AOI22X1 inst_cellmath__37_0_I705 (.Y(N3837), .A0(N3827), .A1(N3983), .B0(N3793), .B1(N3777));
AOI22X1 inst_cellmath__37_0_I706 (.Y(N3882), .A0(N3827), .A1(N3810), .B0(N3841), .B1(N3777));
AOI22XL inst_cellmath__37_0_I707 (.Y(N3929), .A0(N3827), .A1(N3861), .B0(N3885), .B1(N3777));
AOI22XL inst_cellmath__37_0_I708 (.Y(N3979), .A0(N3827), .A1(N3905), .B0(N3777), .B1(N3932));
AOI22XL inst_cellmath__37_0_I709 (.Y(N3807), .A0(N3827), .A1(N3953), .B0(N3777), .B1(N3983));
AOI22X1 inst_cellmath__37_0_I710 (.Y(N3858), .A0(N3827), .A1(N3784), .B0(N3810), .B1(N3777));
AOI22XL inst_cellmath__37_0_I711 (.Y(N3901), .A0(N3827), .A1(N3833), .B0(N3777), .B1(N3861));
AOI22X1 inst_cellmath__37_0_I712 (.Y(N3950), .A0(N3827), .A1(N3876), .B0(N3905), .B1(N3777));
AOI22X1 inst_cellmath__37_0_I713 (.Y(N3781), .A0(N3827), .A1(N3925), .B0(N3953), .B1(N3777));
AOI22X1 inst_cellmath__37_0_I714 (.Y(N3830), .A0(N3827), .A1(N3973), .B0(N3777), .B1(N3784));
AOI22X1 inst_cellmath__37_0_I715 (.Y(N3873), .A0(N3827), .A1(N3803), .B0(N3777), .B1(N3833));
AOI22XL inst_cellmath__37_0_I716 (.Y(N3922), .A0(N3827), .A1(N3852), .B0(N3876), .B1(N3777));
AOI22XL inst_cellmath__37_0_I717 (.Y(N3970), .A0(N3827), .A1(N3897), .B0(N3925), .B1(N3777));
AOI22X1 inst_cellmath__37_0_I718 (.Y(N3800), .A0(N3827), .A1(N3943), .B0(N3777), .B1(N3973));
AOI22X1 inst_cellmath__37_0_I719 (.Y(N3849), .A0(N3827), .A1(N3775), .B0(N3803), .B1(N3777));
AOI22X1 inst_cellmath__37_0_I720 (.Y(N3894), .A0(N3822), .A1(N3827), .B0(N3777), .B1(N3852));
AOI22XL inst_cellmath__37_0_I721 (.Y(N3940), .A0(N3827), .A1(N3868), .B0(N3897), .B1(N3777));
AOI22XL inst_cellmath__37_0_I722 (.Y(N3772), .A0(N3827), .A1(N3947), .B0(N3777), .B1(N3943));
NAND2XL inst_cellmath__37_0_I723 (.Y(N3819), .A(N3775), .B(N3777));
NAND2XL inst_cellmath__37_0_I724 (.Y(N3912), .A(N3822), .B(N3777));
NAND2XL inst_cellmath__37_0_I725 (.Y(N3794), .A(N3868), .B(N3777));
NAND2XL inst_cellmath__37_0_I726 (.Y(N3886), .A(N3947), .B(N3777));
CLKINVX4 inst_cellmath__37_0_I727 (.Y(N3918), .A(inst_cellmath__35[1]));
INVX1 inst_cellmath__37_0_I728 (.Y(N3967), .A(N3918));
NOR2XL inst_cellmath__37_0_I729 (.Y(N3778), .A(N3918), .B(N3966));
NOR2XL inst_cellmath__37_0_I730 (.Y(N3919), .A(N3918), .B(N3845));
AOI22XL inst_cellmath__37_0_I731 (.Y(N3847), .A0(N3918), .A1(N3966), .B0(N3937), .B1(N3967));
AOI22XL inst_cellmath__37_0_I732 (.Y(N3891), .A0(N3918), .A1(N3845), .B0(N3815), .B1(N3967));
AOI22X1 inst_cellmath__37_0_I733 (.Y(N3938), .A0(N3918), .A1(N3937), .B0(N3909), .B1(N3967));
AOI22XL inst_cellmath__37_0_I734 (.Y(N3769), .A0(N3815), .A1(N3918), .B0(N3967), .B1(N3957));
AOI22X1 inst_cellmath__37_0_I735 (.Y(N3817), .A0(N3918), .A1(N3909), .B0(N3967), .B1(N3790));
AOI22XL inst_cellmath__37_0_I736 (.Y(N3865), .A0(N3918), .A1(N3957), .B0(N3837), .B1(N3967));
AOI22X1 inst_cellmath__37_0_I737 (.Y(N3910), .A0(N3918), .A1(N3790), .B0(N3967), .B1(N3882));
AOI22XL inst_cellmath__37_0_I738 (.Y(N3958), .A0(N3918), .A1(N3837), .B0(N3967), .B1(N3929));
AOI22XL inst_cellmath__37_0_I739 (.Y(N3792), .A0(N3918), .A1(N3882), .B0(N3967), .B1(N3979));
AOI22XL inst_cellmath__37_0_I740 (.Y(N3839), .A0(N3918), .A1(N3929), .B0(N3807), .B1(N3967));
AOI22X1 inst_cellmath__37_0_I741 (.Y(N3884), .A0(N3918), .A1(N3979), .B0(N3967), .B1(N3858));
AOI22X1 inst_cellmath__37_0_I742 (.Y(N3931), .A0(N3807), .A1(N3918), .B0(N3967), .B1(N3901));
AOI22XL inst_cellmath__37_0_I743 (.Y(N3982), .A0(N3918), .A1(N3858), .B0(N3950), .B1(N3967));
AOI22XL inst_cellmath__37_0_I744 (.Y(N3809), .A0(N3918), .A1(N3901), .B0(N3781), .B1(N3967));
AOI22X1 inst_cellmath__37_0_I745 (.Y(N3860), .A0(N3918), .A1(N3950), .B0(N3967), .B1(N3830));
AOI22X1 inst_cellmath__37_0_I746 (.Y(N3903), .A0(N3918), .A1(N3781), .B0(N3967), .B1(N3873));
AOI22XL inst_cellmath__37_0_I747 (.Y(N3952), .A0(N3918), .A1(N3830), .B0(N3967), .B1(N3922));
AOI22XL inst_cellmath__37_0_I748 (.Y(N3783), .A0(N3918), .A1(N3873), .B0(N3967), .B1(N3970));
AOI22X1 inst_cellmath__37_0_I749 (.Y(N3832), .A0(N3918), .A1(N3922), .B0(N3800), .B1(N3967));
AOI22X1 inst_cellmath__37_0_I750 (.Y(N3875), .A0(N3918), .A1(N3970), .B0(N3967), .B1(N3849));
AOI22X1 inst_cellmath__37_0_I751 (.Y(N3924), .A0(N3918), .A1(N3800), .B0(N3967), .B1(N3894));
AOI22X1 inst_cellmath__37_0_I752 (.Y(N3972), .A0(N3918), .A1(N3849), .B0(N3967), .B1(N3940));
AOI22X1 inst_cellmath__37_0_I753 (.Y(N3802), .A0(N3918), .A1(N3894), .B0(N3772), .B1(N3967));
AOI22X1 inst_cellmath__37_0_I754 (.Y(N3851), .A0(N3918), .A1(N3940), .B0(N3819), .B1(N3967));
AOI22XL inst_cellmath__37_0_I755 (.Y(N3896), .A0(N3918), .A1(N3772), .B0(N3912), .B1(N3967));
AOI22XL inst_cellmath__37_0_I756 (.Y(N3942), .A0(N3918), .A1(N3819), .B0(N3794), .B1(N3967));
AOI22XL inst_cellmath__37_0_I757 (.Y(N3774), .A0(N3918), .A1(N3912), .B0(N3886), .B1(N3967));
NOR2XL inst_cellmath__37_0_I758 (.Y(N3821), .A(N3967), .B(N3794));
NOR2XL inst_cellmath__37_0_I759 (.Y(N3963), .A(N3967), .B(N3886));
CLKINVX4 inst_cellmath__37_0_I760 (.Y(N3846), .A(inst_cellmath__35[4]));
CLKINVX4 inst_cellmath__37_0_I761 (.Y(N3890), .A(N3846));
NAND2XL inst_cellmath__37_0_I762 (.Y(N3961), .A(N3890), .B(N3778));
NAND2XL inst_cellmath__37_0_I763 (.Y(N3842), .A(N3890), .B(N3919));
NAND2XL inst_cellmath__37_0_I764 (.Y(N3934), .A(N3890), .B(N3847));
NAND2XL inst_cellmath__37_0_I765 (.Y(N3812), .A(N3890), .B(N3891));
NAND2XL inst_cellmath__37_0_I766 (.Y(N3906), .A(N3890), .B(N3938));
NAND2XL inst_cellmath__37_0_I767 (.Y(N3786), .A(N3890), .B(N3769));
NAND2XL inst_cellmath__37_0_I768 (.Y(N3878), .A(N3890), .B(N3817));
NAND2X1 inst_cellmath__37_0_I769 (.Y(N3975), .A(N3890), .B(N3865));
NAND2X1 inst_cellmath__37_0_I770 (.Y(N3854), .A(N3890), .B(N3910));
NAND2XL inst_cellmath__37_0_I771 (.Y(N3945), .A(N3890), .B(N3958));
NAND2X1 inst_cellmath__37_0_I772 (.Y(N3825), .A(N3890), .B(N3792));
NAND2X1 inst_cellmath__37_0_I773 (.Y(N3916), .A(N3890), .B(N3839));
NAND2X1 inst_cellmath__37_0_I774 (.Y(N3795), .A(N3890), .B(N3884));
NAND2X1 inst_cellmath__37_0_I775 (.Y(N3888), .A(N3890), .B(N3931));
NAND2X1 inst_cellmath__37_0_I776 (.Y(N3766), .A(N3890), .B(N3982));
NAND2XL inst_cellmath__37_0_I777 (.Y(N3863), .A(N3890), .B(N3809));
AOI22X1 inst_cellmath__37_0_I778 (.Y(N3955), .A0(N3890), .A1(N3860), .B0(N3778), .B1(N3846));
AOI22X1 inst_cellmath__37_0_I779 (.Y(N3788), .A0(N3890), .A1(N3903), .B0(N3919), .B1(N3846));
AOI22X1 inst_cellmath__37_0_I780 (.Y(N3835), .A0(N3890), .A1(N3952), .B0(N3846), .B1(N3847));
AOI22X1 inst_cellmath__37_0_I781 (.Y(N3880), .A0(N3890), .A1(N3783), .B0(N3846), .B1(N3891));
AOI22X2 inst_cellmath__37_0_I782 (.Y(N3927), .A0(N3890), .A1(N3832), .B0(N3846), .B1(N3938));
AOI22X1 inst_cellmath__37_0_I783 (.Y(N3977), .A0(N3890), .A1(N3875), .B0(N3846), .B1(N3769));
AOI22X1 inst_cellmath__37_0_I784 (.Y(N3805), .A0(N3890), .A1(N3924), .B0(N3846), .B1(N3817));
AOI22XL inst_cellmath__37_0_I785 (.Y(N3856), .A0(N3890), .A1(N3972), .B0(N3846), .B1(N3865));
AOI22X1 inst_cellmath__37_0_I786 (.Y(N3899), .A0(N3890), .A1(N3802), .B0(N3846), .B1(N3910));
AOI22XL inst_cellmath__37_0_I787 (.Y(N3948), .A0(N3851), .A1(N3890), .B0(N3846), .B1(N3958));
AOI22XL inst_cellmath__37_0_I788 (.Y(N3779), .A0(N3896), .A1(N3890), .B0(N3846), .B1(N3792));
AOI22XL inst_cellmath__37_0_I789 (.Y(N3828), .A0(N3942), .A1(N3890), .B0(N3846), .B1(N3839));
AOI22XL inst_cellmath__37_0_I790 (.Y(N3871), .A0(N3774), .A1(N3890), .B0(N3846), .B1(N3884));
AOI22XL inst_cellmath__37_0_I791 (.Y(N3920), .A0(N3890), .A1(N3821), .B0(N3931), .B1(N3846));
AOI22XL inst_cellmath__37_0_I792 (.Y(N3968), .A0(N3963), .A1(N3890), .B0(N3846), .B1(N3982));
NAND2XL inst_cellmath__37_0_I793 (.Y(N3798), .A(N3846), .B(N3809));
NAND2XL inst_cellmath__37_0_I794 (.Y(N3892), .A(N3860), .B(N3846));
NAND2XL inst_cellmath__37_0_I795 (.Y(N3770), .A(N3903), .B(N3846));
NAND2XL inst_cellmath__37_0_I796 (.Y(N3866), .A(N3846), .B(N3952));
NAND2XL inst_cellmath__37_0_I797 (.Y(N3960), .A(N3846), .B(N3783));
NAND2XL inst_cellmath__37_0_I798 (.Y(N3840), .A(N3846), .B(N3832));
NAND2XL inst_cellmath__37_0_I799 (.Y(N3933), .A(N3875), .B(N3846));
NAND2XL inst_cellmath__37_0_I800 (.Y(N3811), .A(N3924), .B(N3846));
NAND2XL inst_cellmath__37_0_I801 (.Y(N3904), .A(N3972), .B(N3846));
NAND2XL inst_cellmath__37_0_I802 (.Y(N3785), .A(N3846), .B(N3802));
NAND2XL inst_cellmath__37_0_I803 (.Y(N3877), .A(N3851), .B(N3846));
NAND2XL inst_cellmath__37_0_I804 (.Y(N3974), .A(N3896), .B(N3846));
NAND2XL inst_cellmath__37_0_I805 (.Y(N3853), .A(N3942), .B(N3846));
NAND2XL inst_cellmath__37_0_I806 (.Y(N3944), .A(N3774), .B(N3846));
NAND2XL inst_cellmath__37_0_I807 (.Y(N3823), .A(N3821), .B(N3846));
NAND2XL inst_cellmath__37_0_I808 (.Y(N3914), .A(N3963), .B(N3846));
CLKINVX6 inst_cellmath__37_0_I2643 (.Y(N3768), .A(inst_cellmath__35[3]));
INVX1 inst_cellmath__37_0_I811 (.Y(N3816), .A(N3768));
NOR2XL inst_cellmath__37_0_I812 (.Y(inst_cellmath__37[0]), .A(N3768), .B(N3786));
NOR2X1 inst_cellmath__37_0_I813 (.Y(inst_cellmath__37[1]), .A(N3768), .B(N3878));
NOR2X1 inst_cellmath__37_0_I814 (.Y(inst_cellmath__37[2]), .A(N3768), .B(N3975));
AOI22XL inst_cellmath__37_0_I815 (.Y(inst_cellmath__37[3]), .A0(N3961), .A1(N3768), .B0(N3816), .B1(N3854));
AOI22XL inst_cellmath__37_0_I816 (.Y(inst_cellmath__37[4]), .A0(N3768), .A1(N3842), .B0(N3945), .B1(N3816));
AOI22X1 inst_cellmath__37_0_I817 (.Y(inst_cellmath__37[5]), .A0(N3768), .A1(N3934), .B0(N3816), .B1(N3825));
AOI22X1 inst_cellmath__37_0_I818 (.Y(inst_cellmath__37[6]), .A0(N3768), .A1(N3812), .B0(N3816), .B1(N3916));
AOI22X1 inst_cellmath__37_0_I819 (.Y(inst_cellmath__37[7]), .A0(N3768), .A1(N3906), .B0(N3816), .B1(N3795));
AOI22XL inst_cellmath__37_0_I820 (.Y(inst_cellmath__37[8]), .A0(N3768), .A1(N3786), .B0(N3816), .B1(N3888));
AOI22X1 inst_cellmath__37_0_I821 (.Y(inst_cellmath__37[9]), .A0(N3768), .A1(N3878), .B0(N3816), .B1(N3766));
AOI22X1 inst_cellmath__37_0_I822 (.Y(inst_cellmath__37[10]), .A0(N3768), .A1(N3975), .B0(N3816), .B1(N3863));
AOI22X1 inst_cellmath__37_0_I824 (.Y(inst_cellmath__37[12]), .A0(N3768), .A1(N3945), .B0(N3816), .B1(N3788));
AOI22X1 inst_cellmath__37_0_I829 (.Y(inst_cellmath__37[17]), .A0(N3768), .A1(N3766), .B0(N3816), .B1(N3805));
AOI22X1 inst_cellmath__37_0_I831 (.Y(inst_cellmath__37[19]), .A0(N3768), .A1(N3955), .B0(N3816), .B1(N3899));
AOI22XL inst_cellmath__37_0_I836 (.Y(inst_cellmath__37[24]), .A0(N3768), .A1(N3977), .B0(N3920), .B1(N3816));
AOI22XL inst_cellmath__37_0_I837 (.Y(inst_cellmath__37[25]), .A0(N3768), .A1(N3805), .B0(N3968), .B1(N3816));
AOI22XL inst_cellmath__37_0_I838 (.Y(inst_cellmath__37[26]), .A0(N3768), .A1(N3856), .B0(N3798), .B1(N3816));
AOI22XL inst_cellmath__37_0_I839 (.Y(inst_cellmath__37[27]), .A0(N3768), .A1(N3899), .B0(N3892), .B1(N3816));
AOI22XL inst_cellmath__37_0_I840 (.Y(inst_cellmath__37[28]), .A0(N3768), .A1(N3948), .B0(N3770), .B1(N3816));
AOI22XL inst_cellmath__37_0_I841 (.Y(inst_cellmath__37[29]), .A0(N3768), .A1(N3779), .B0(N3866), .B1(N3816));
AOI22XL inst_cellmath__37_0_I842 (.Y(inst_cellmath__37[30]), .A0(N3768), .A1(N3828), .B0(N3960), .B1(N3816));
AOI22XL inst_cellmath__37_0_I843 (.Y(inst_cellmath__37[31]), .A0(N3768), .A1(N3871), .B0(N3840), .B1(N3816));
AOI22XL inst_cellmath__37_0_I844 (.Y(inst_cellmath__37[32]), .A0(N3768), .A1(N3920), .B0(N3933), .B1(N3816));
AOI22XL inst_cellmath__37_0_I845 (.Y(inst_cellmath__37[33]), .A0(N3768), .A1(N3968), .B0(N3811), .B1(N3816));
AOI22XL inst_cellmath__37_0_I846 (.Y(inst_cellmath__37[34]), .A0(N3768), .A1(N3798), .B0(N3904), .B1(N3816));
AOI22XL inst_cellmath__37_0_I847 (.Y(inst_cellmath__37[35]), .A0(N3768), .A1(N3892), .B0(N3785), .B1(N3816));
AOI22XL inst_cellmath__37_0_I848 (.Y(inst_cellmath__37[36]), .A0(N3768), .A1(N3770), .B0(N3877), .B1(N3816));
AOI22XL inst_cellmath__37_0_I849 (.Y(inst_cellmath__37[37]), .A0(N3768), .A1(N3866), .B0(N3974), .B1(N3816));
AOI22XL inst_cellmath__37_0_I850 (.Y(inst_cellmath__37[38]), .A0(N3768), .A1(N3960), .B0(N3853), .B1(N3816));
AOI22XL inst_cellmath__37_0_I851 (.Y(inst_cellmath__37[39]), .A0(N3768), .A1(N3840), .B0(N3944), .B1(N3816));
AOI22XL inst_cellmath__37_0_I852 (.Y(inst_cellmath__37[40]), .A0(N3768), .A1(N3933), .B0(N3823), .B1(N3816));
AOI22XL inst_cellmath__37_0_I853 (.Y(inst_cellmath__37[41]), .A0(N3768), .A1(N3811), .B0(N3914), .B1(N3816));
OR2X1 cynw_cm_float_add2_ieee_I6905 (.Y(inst_cellmath__31), .A(inst_cellmath__11), .B(inst_cellmath__16));
NOR2X1 inst_cellmath__33_49_24_I2644 (.Y(N4205), .A(inst_cellmath__31), .B(inst_cellmath__30));
AND2XL inst_cellmath__33_49_24_I863 (.Y(inst_cellmath__33[24]), .A(N4205), .B(inst_cellmath__37[24]));
AND2XL inst_cellmath__33_49_24_I864 (.Y(inst_cellmath__33[25]), .A(N4205), .B(inst_cellmath__37[25]));
AND2XL inst_cellmath__33_49_24_I865 (.Y(inst_cellmath__33[26]), .A(N4205), .B(inst_cellmath__37[26]));
AND2XL inst_cellmath__33_49_24_I866 (.Y(inst_cellmath__33[27]), .A(N4205), .B(inst_cellmath__37[27]));
AND2XL inst_cellmath__33_49_24_I867 (.Y(inst_cellmath__33[28]), .A(N4205), .B(inst_cellmath__37[28]));
AND2XL inst_cellmath__33_49_24_I869 (.Y(inst_cellmath__33[30]), .A(N4205), .B(inst_cellmath__37[30]));
AND2XL inst_cellmath__33_49_24_I871 (.Y(inst_cellmath__33[32]), .A(N4205), .B(inst_cellmath__37[32]));
AND2XL inst_cellmath__33_49_24_I873 (.Y(inst_cellmath__33[34]), .A(N4205), .B(inst_cellmath__37[34]));
AND2XL inst_cellmath__33_49_24_I875 (.Y(inst_cellmath__33[36]), .A(N4205), .B(inst_cellmath__37[36]));
AND2XL inst_cellmath__33_49_24_I877 (.Y(inst_cellmath__33[38]), .A(N4205), .B(inst_cellmath__37[38]));
AND2XL inst_cellmath__33_49_24_I879 (.Y(inst_cellmath__33[40]), .A(N4205), .B(inst_cellmath__37[40]));
AND2XL inst_cellmath__33_49_24_I880 (.Y(inst_cellmath__33[41]), .A(N4205), .B(inst_cellmath__37[41]));
NOR3BXL inst_cellmath__33_49_24_I2645 (.Y(inst_cellmath__33[42]), .AN(N4205), .B(N3816), .C(N3904));
NOR3BXL inst_cellmath__33_49_24_I2646 (.Y(inst_cellmath__33[43]), .AN(N4205), .B(N3816), .C(N3785));
NOR3BXL inst_cellmath__33_49_24_I2647 (.Y(inst_cellmath__33[44]), .AN(N4205), .B(N3816), .C(N3877));
NOR3BXL inst_cellmath__33_49_24_I2648 (.Y(inst_cellmath__33[45]), .AN(N4205), .B(N3816), .C(N3974));
NOR3BXL inst_cellmath__33_49_24_I2649 (.Y(inst_cellmath__33[46]), .AN(N4205), .B(N3816), .C(N3853));
NOR3BXL inst_cellmath__33_49_24_I2650 (.Y(inst_cellmath__33[47]), .AN(N4205), .B(N3816), .C(N3944));
NOR3BXL inst_cellmath__33_49_24_I2651 (.Y(inst_cellmath__33[48]), .AN(N4205), .B(N3816), .C(N3823));
NOR3BXL inst_cellmath__33_49_24_I2652 (.Y(inst_cellmath__33[49]), .AN(N4205), .B(N3816), .C(N3914));
NOR2X1 inst_cellmath__42__22__I889 (.Y(N4261), .A(inst_cellmath__30), .B(inst_cellmath__37[0]));
NOR2X2 inst_cellmath__42__22__I890 (.Y(N4271), .A(inst_cellmath__37[1]), .B(inst_cellmath__37[2]));
NAND2X2 inst_cellmath__42__22__I891 (.Y(N4282), .A(N4261), .B(N4271));
NOR2X1 inst_cellmath__42__22__I892 (.Y(N4291), .A(inst_cellmath__37[3]), .B(inst_cellmath__37[7]));
NOR2X1 inst_cellmath__42__22__I893 (.Y(N4300), .A(inst_cellmath__37[9]), .B(inst_cellmath__37[5]));
NOR2X1 inst_cellmath__42__22__I894 (.Y(N4265), .A(inst_cellmath__37[6]), .B(inst_cellmath__37[8]));
NOR2X1 inst_cellmath__42__22__I895 (.Y(N4274), .A(inst_cellmath__37[4]), .B(inst_cellmath__37[10]));
NOR2X1 inst_cellmath__42__22__I896 (.Y(N4294), .A(inst_cellmath__37[12]), .B(inst_cellmath__37[17]));
NOR2X2 inst_cellmath__42__22__I897 (.Y(N4279), .A(N4282), .B(inst_cellmath__37[19]));
AOI22XL cynw_cm_float_add2_ieee_I6906 (.Y(N12033), .A0(N3768), .A1(N3854), .B0(N3955), .B1(N3816));
AOI22X1 cynw_cm_float_add2_ieee_I6907 (.Y(N12046), .A0(N3768), .A1(N3825), .B0(N3816), .B1(N3835));
AOI22X1 cynw_cm_float_add2_ieee_I6908 (.Y(N12060), .A0(N3768), .A1(N3916), .B0(N3816), .B1(N3880));
AOI22X2 cynw_cm_float_add2_ieee_I6909 (.Y(N12073), .A0(N3768), .A1(N3795), .B0(N3816), .B1(N3927));
AOI22X1 cynw_cm_float_add2_ieee_I6910 (.Y(N12086), .A0(N3768), .A1(N3888), .B0(N3816), .B1(N3977));
AOI22XL cynw_cm_float_add2_ieee_I6911 (.Y(N12038), .A0(N3768), .A1(N3863), .B0(N3816), .B1(N3856));
AOI22X1 cynw_cm_float_add2_ieee_I6912 (.Y(N12052), .A0(N3768), .A1(N3788), .B0(N3948), .B1(N3816));
AOI22X2 cynw_cm_float_add2_ieee_I6913 (.Y(N12066), .A0(N3835), .A1(N3768), .B0(N3816), .B1(N3779));
AOI22X1 cynw_cm_float_add2_ieee_I6914 (.Y(N12079), .A0(N3768), .A1(N3880), .B0(N3816), .B1(N3828));
AOI22X1 cynw_cm_float_add2_ieee_I6915 (.Y(N12092), .A0(N3768), .A1(N3927), .B0(N3816), .B1(N3871));
NAND2X1 cynw_cm_float_add2_ieee_I6916 (.Y(N12043), .A(N4291), .B(N4300));
NAND2X1 cynw_cm_float_add2_ieee_I6917 (.Y(N12057), .A(N4265), .B(N4274));
NAND2X2 cynw_cm_float_add2_ieee_I6918 (.Y(N12070), .A(N4294), .B(N4279));
NOR4X2 cynw_cm_float_add2_ieee_I6919 (.Y(N12083), .A(N12073), .B(N12086), .C(N12033), .D(N12046));
NOR3X2 cynw_cm_float_add2_ieee_I6920 (.Y(N12036), .A(N12038), .B(N12060), .C(N12043));
NOR3X2 cynw_cm_float_add2_ieee_I6921 (.Y(N12049), .A(N12092), .B(N12079), .C(N12057));
NOR3X4 cynw_cm_float_add2_ieee_I6922 (.Y(N12063), .A(N12052), .B(N12066), .C(N12070));
NAND2X2 cynw_cm_float_add2_ieee_I6923 (.Y(N12076), .A(N12036), .B(N12083));
NAND2X4 cynw_cm_float_add2_ieee_I6924 (.Y(N12088), .A(N12049), .B(N12063));
NOR2X4 cynw_cm_float_add2_ieee_I6925 (.Y(N12091), .A(N12076), .B(N12088));
INVXL cynw_cm_float_add2_ieee_I7115 (.Y(N12585), .A(rm[2]));
INVXL cynw_cm_float_add2_ieee_I7116 (.Y(N12547), .A(rm[1]));
NOR3BXL cynw_cm_float_add2_ieee_I7117 (.Y(inst_cellmath__6), .AN(N12585), .B(N12547), .C(rm[0]));
INVXL buf1_A_I7321 (.Y(N12695), .A(inst_cellmath__32));
INVXL buf1_A_I7322 (.Y(N12595), .A(N12695));
INVXL cynw_cm_float_add2_ieee_I7121 (.Y(N12582), .A(N12595));
NOR2BX1 cynw_cm_float_add2_ieee_I7211 (.Y(N12548), .AN(a_sign), .B(N12582));
AND2XL cynw_cm_float_add2_ieee_I7123 (.Y(N12565), .A(b_sign), .B(N12582));
MX2XL cynw_cm_float_add2_ieee_I7124 (.Y(inst_cellmath__48), .A(a_sign), .B(b_sign), .S0(N12582));
MX2XL cynw_cm_float_add2_ieee_I918 (.Y(N660), .A(a_man[5]), .B(b_man[5]), .S0(N3695));
INVX1 inst_cellmath__44_0_I909 (.Y(N4328), .A(inst_cellmath__39[25]));
NAND2XL node_cs_const1_cs_ii_A_I7323 (.Y(N12699), .A(N4205), .B(inst_cellmath__37[31]));
XOR2XL node_cs_const1_cs_ii_A_I7324 (.Y(inst_cellmath__39[6]), .A(N4328), .B(N12699));
XNOR2X1 inst_cellmath__45_0_I968 (.Y(N4511), .A(inst_cellmath__39[6]), .B(N660));
MX2XL cynw_cm_float_add2_ieee_I917 (.Y(N659), .A(a_man[4]), .B(b_man[4]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I942 (.Y(inst_cellmath__39[5]), .A(N4328), .B(inst_cellmath__33[30]));
MX2XL cynw_cm_float_add2_ieee_I916 (.Y(N658), .A(a_man[3]), .B(b_man[3]), .S0(N3695));
NAND2XL node_cs_const1_cs_ii_A_I7325 (.Y(N12706), .A(N4205), .B(inst_cellmath__37[29]));
XOR2XL node_cs_const1_cs_ii_A_I7326 (.Y(inst_cellmath__39[4]), .A(N4328), .B(N12706));
XNOR2X1 inst_cellmath__45_0_I966 (.Y(N4524), .A(inst_cellmath__39[4]), .B(N658));
MX2XL cynw_cm_float_add2_ieee_I915 (.Y(N657), .A(a_man[2]), .B(b_man[2]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I940 (.Y(inst_cellmath__39[3]), .A(N4328), .B(inst_cellmath__33[28]));
MX2XL cynw_cm_float_add2_ieee_I914 (.Y(N656), .A(a_man[1]), .B(b_man[1]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I939 (.Y(inst_cellmath__39[2]), .A(N4328), .B(inst_cellmath__33[27]));
XNOR2X1 inst_cellmath__45_0_I964 (.Y(N4541), .A(inst_cellmath__39[2]), .B(N656));
MX2XL cynw_cm_float_add2_ieee_I913 (.Y(N655), .A(N11653), .B(b_man[0]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I938 (.Y(inst_cellmath__39[1]), .A(N4328), .B(inst_cellmath__33[26]));
XNOR2X1 inst_cellmath__39__19__2mx_I937 (.Y(inst_cellmath__39[0]), .A(inst_cellmath__33[25]), .B(N4328));
NOR2X6 cynw_cm_float_add2_ieee_I7139 (.Y(inst_cellmath__42), .A(inst_cellmath__31), .B(N12091));
NOR3X8 inst_cellmath__44_0_I910 (.Y(inst_cellmath__44), .A(N4328), .B(inst_cellmath__33[24]), .C(inst_cellmath__42));
NAND2X6 inst_cellmath__45_0_I962 (.Y(N4556), .A(inst_cellmath__39[0]), .B(inst_cellmath__44));
CLKXOR2X2 inst_cellmath__45_0_I963 (.Y(N4618), .A(N655), .B(inst_cellmath__39[1]));
AOI2BB2X4 inst_cellmath__45_0_I990 (.Y(N4575), .A0N(inst_cellmath__39[1]), .A1N(N655), .B0(N4556), .B1(N4618));
OAI22X4 inst_cellmath__45_0_I991 (.Y(N4540), .A0(N4541), .A1(N4575), .B0(inst_cellmath__39[2]), .B1(N656));
CLKXOR2X2 inst_cellmath__45_0_I965 (.Y(N4601), .A(N657), .B(inst_cellmath__39[3]));
AOI2BB2X4 inst_cellmath__45_0_I992 (.Y(N4510), .A0N(inst_cellmath__39[3]), .A1N(N657), .B0(N4540), .B1(N4601));
OAI22X4 inst_cellmath__45_0_I993 (.Y(N4592), .A0(N4524), .A1(N4510), .B0(inst_cellmath__39[4]), .B1(N658));
CLKXOR2X2 inst_cellmath__45_0_I967 (.Y(N4582), .A(N659), .B(inst_cellmath__39[5]));
AOI2BB2X4 inst_cellmath__45_0_I994 (.Y(N4537), .A0N(inst_cellmath__39[5]), .A1N(N659), .B0(N4592), .B1(N4582));
OAI22X4 inst_cellmath__45_0_I995 (.Y(N4604), .A0(N4511), .A1(N4537), .B0(inst_cellmath__39[6]), .B1(N660));
MX2XL cynw_cm_float_add2_ieee_I919 (.Y(N661), .A(a_man[6]), .B(b_man[6]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I944 (.Y(inst_cellmath__39[7]), .A(inst_cellmath__33[32]), .B(N4328));
CLKXOR2X2 inst_cellmath__45_0_I969 (.Y(N4566), .A(N661), .B(inst_cellmath__39[7]));
XNOR2X1 inst_cellmath__45_0_I1020 (.Y(inst_cellmath__45[7]), .A(N4604), .B(N4566));
XNOR2X1 inst_cellmath__45_0_I1019 (.Y(inst_cellmath__45[6]), .A(N4537), .B(N4511));
NOR2XL inst_cellmath__49_0_I1050 (.Y(N4752), .A(inst_cellmath__45[7]), .B(inst_cellmath__45[6]));
XNOR2X1 inst_cellmath__45_0_I1016 (.Y(inst_cellmath__45[3]), .A(N4540), .B(N4601));
XNOR2X1 inst_cellmath__45_0_I1015 (.Y(inst_cellmath__45[2]), .A(N4575), .B(N4541));
NOR2XL inst_cellmath__49_0_I1045 (.Y(N4725), .A(inst_cellmath__45[3]), .B(inst_cellmath__45[2]));
XNOR2X1 inst_cellmath__45_0_I1018 (.Y(inst_cellmath__45[5]), .A(N4592), .B(N4582));
XNOR2X1 inst_cellmath__45_0_I1017 (.Y(inst_cellmath__45[4]), .A(N4510), .B(N4524));
NOR2XL inst_cellmath__49_0_I1046 (.Y(N4744), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[4]));
NAND2BXL inst_cellmath__49_0_I1072 (.Y(N4792), .AN(N4725), .B(N4744));
MX2XL cynw_cm_float_add2_ieee_I920 (.Y(N662), .A(a_man[7]), .B(b_man[7]), .S0(N3695));
NAND2XL node_cs_const1_cs_ii_A_I7327 (.Y(N12713), .A(N4205), .B(inst_cellmath__37[33]));
XOR2XL node_cs_const1_cs_ii_A_I7328 (.Y(inst_cellmath__39[8]), .A(N4328), .B(N12713));
XNOR2X1 inst_cellmath__45_0_I970 (.Y(N4623), .A(inst_cellmath__39[8]), .B(N662));
AOI2BB2X4 inst_cellmath__45_0_I996 (.Y(N4534), .A0N(N661), .A1N(inst_cellmath__39[7]), .B0(N4604), .B1(N4566));
OAI22X4 inst_cellmath__45_0_I997 (.Y(N4585), .A0(N4623), .A1(N4534), .B0(inst_cellmath__39[8]), .B1(N662));
MX2XL cynw_cm_float_add2_ieee_I921 (.Y(N663), .A(a_man[8]), .B(b_man[8]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I946 (.Y(inst_cellmath__39[9]), .A(inst_cellmath__33[34]), .B(N4328));
CLKXOR2X2 inst_cellmath__45_0_I971 (.Y(N4546), .A(N663), .B(inst_cellmath__39[9]));
XNOR2X1 inst_cellmath__45_0_I1022 (.Y(inst_cellmath__45[9]), .A(N4585), .B(N4546));
XNOR2X1 inst_cellmath__45_0_I1021 (.Y(inst_cellmath__45[8]), .A(N4534), .B(N4623));
NOR2XL inst_cellmath__49_0_I1051 (.Y(N4771), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[8]));
OAI2BB1X1 inst_cellmath__49_0_I1100 (.Y(N4784), .A0N(N4752), .A1N(N4792), .B0(N4771));
MX2XL cynw_cm_float_add2_ieee_I928 (.Y(N670), .A(a_man[15]), .B(b_man[15]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I953 (.Y(inst_cellmath__39[16]), .A(inst_cellmath__33[41]), .B(N4328));
XNOR2X1 inst_cellmath__45_0_I978 (.Y(N4554), .A(N670), .B(inst_cellmath__39[16]));
MX2XL cynw_cm_float_add2_ieee_I927 (.Y(N669), .A(a_man[14]), .B(b_man[14]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I952 (.Y(inst_cellmath__39[15]), .A(inst_cellmath__33[40]), .B(N4328));
MX2XL cynw_cm_float_add2_ieee_I926 (.Y(N668), .A(a_man[13]), .B(b_man[13]), .S0(N3695));
NAND2XL node_cs_const1_cs_ii_A_I7329 (.Y(N12720), .A(N4205), .B(inst_cellmath__37[39]));
XOR2XL node_cs_const1_cs_ii_A_I7330 (.Y(inst_cellmath__39[14]), .A(N4328), .B(N12720));
XNOR2X1 inst_cellmath__45_0_I976 (.Y(N4572), .A(inst_cellmath__39[14]), .B(N668));
MX2XL cynw_cm_float_add2_ieee_I925 (.Y(N667), .A(a_man[12]), .B(b_man[12]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I950 (.Y(inst_cellmath__39[13]), .A(N4328), .B(inst_cellmath__33[38]));
MX2XL cynw_cm_float_add2_ieee_I924 (.Y(N666), .A(a_man[11]), .B(b_man[11]), .S0(N3695));
NAND2XL node_cs_const1_cs_ii_A_I7331 (.Y(N12727), .A(N4205), .B(inst_cellmath__37[37]));
XOR2XL node_cs_const1_cs_ii_A_I7332 (.Y(inst_cellmath__39[12]), .A(N4328), .B(N12727));
XNOR2X1 inst_cellmath__45_0_I974 (.Y(N4594), .A(inst_cellmath__39[12]), .B(N666));
MX2XL cynw_cm_float_add2_ieee_I923 (.Y(N665), .A(a_man[10]), .B(b_man[10]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I948 (.Y(inst_cellmath__39[11]), .A(N4328), .B(inst_cellmath__33[36]));
MX2XL cynw_cm_float_add2_ieee_I922 (.Y(N664), .A(a_man[9]), .B(b_man[9]), .S0(N3695));
NAND2XL node_cs_const1_cs_ii_A_I7333 (.Y(N12734), .A(N4205), .B(inst_cellmath__37[35]));
XOR2XL node_cs_const1_cs_ii_A_I7334 (.Y(inst_cellmath__39[10]), .A(N4328), .B(N12734));
XNOR2X1 inst_cellmath__45_0_I972 (.Y(N4609), .A(inst_cellmath__39[10]), .B(N664));
AOI2BB2X4 inst_cellmath__45_0_I998 (.Y(N4631), .A0N(inst_cellmath__39[9]), .A1N(N663), .B0(N4585), .B1(N4546));
OAI22X4 inst_cellmath__45_0_I999 (.Y(N4529), .A0(N4609), .A1(N4631), .B0(inst_cellmath__39[10]), .B1(N664));
CLKXOR2X2 inst_cellmath__45_0_I973 (.Y(N4530), .A(N665), .B(inst_cellmath__39[11]));
AOI2BB2X4 inst_cellmath__45_0_I1000 (.Y(N4561), .A0N(inst_cellmath__39[11]), .A1N(N665), .B0(N4529), .B1(N4530));
OAI22X4 inst_cellmath__45_0_I1001 (.Y(N4576), .A0(N4594), .A1(N4561), .B0(inst_cellmath__39[12]), .B1(N666));
CLKXOR2X2 inst_cellmath__45_0_I975 (.Y(N4518), .A(N667), .B(inst_cellmath__39[13]));
AOI2BB2X4 inst_cellmath__45_0_I1002 (.Y(N4593), .A0N(inst_cellmath__39[13]), .A1N(N667), .B0(N4576), .B1(N4518));
OAI22X4 inst_cellmath__45_0_I1003 (.Y(N4589), .A0(N4572), .A1(N4593), .B0(inst_cellmath__39[14]), .B1(N668));
CLKXOR2X2 inst_cellmath__45_0_I977 (.Y(N4630), .A(N669), .B(inst_cellmath__39[15]));
AOI2BB2X4 inst_cellmath__45_0_I1004 (.Y(N4586), .A0N(inst_cellmath__39[15]), .A1N(N669), .B0(N4589), .B1(N4630));
OAI22X4 inst_cellmath__45_0_I1005 (.Y(N4564), .A0(N4554), .A1(N4586), .B0(inst_cellmath__39[16]), .B1(N670));
MX2XL cynw_cm_float_add2_ieee_I929 (.Y(N671), .A(a_man[16]), .B(b_man[16]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I954 (.Y(inst_cellmath__39[17]), .A(inst_cellmath__33[42]), .B(N4328));
XOR2XL inst_cellmath__45_0_I980 (.Y(N4614), .A(N671), .B(inst_cellmath__39[17]));
XNOR2X1 inst_cellmath__45_0_I1030 (.Y(inst_cellmath__45[17]), .A(N4564), .B(N4614));
XNOR2X1 inst_cellmath__45_0_I1029 (.Y(inst_cellmath__45[16]), .A(N4586), .B(N4554));
NOR2XL inst_cellmath__49_0_I1061 (.Y(N4738), .A(inst_cellmath__45[17]), .B(inst_cellmath__45[16]));
XNOR2X1 inst_cellmath__45_0_I1028 (.Y(inst_cellmath__45[15]), .A(N4589), .B(N4630));
XNOR2X1 inst_cellmath__45_0_I1027 (.Y(inst_cellmath__45[14]), .A(N4593), .B(N4572));
NOR2XL inst_cellmath__49_0_I1060 (.Y(N4717), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[14]));
NAND2XL inst_cellmath__49_0_I1079 (.Y(N4714), .A(N4738), .B(N4717));
XNOR2X1 inst_cellmath__45_0_I1026 (.Y(inst_cellmath__45[13]), .A(N4576), .B(N4518));
XNOR2X1 inst_cellmath__45_0_I1025 (.Y(inst_cellmath__45[12]), .A(N4561), .B(N4594));
NOR2XL inst_cellmath__49_0_I1056 (.Y(N4802), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[12]));
XNOR2X1 inst_cellmath__45_0_I1024 (.Y(inst_cellmath__45[11]), .A(N4529), .B(N4530));
XNOR2X1 inst_cellmath__45_0_I1023 (.Y(inst_cellmath__45[10]), .A(N4631), .B(N4609));
NOR2XL inst_cellmath__49_0_I1055 (.Y(N4782), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[10]));
NAND2XL inst_cellmath__49_0_I1078 (.Y(N4788), .A(N4802), .B(N4782));
NOR2XL inst_cellmath__49_0_I1090 (.Y(N4730), .A(N4714), .B(N4788));
XNOR2X1 inst_cellmath__39__19__2mx_I961 (.Y(inst_cellmath__39[24]), .A(inst_cellmath__33[49]), .B(N4328));
MX2XL cynw_cm_float_add2_ieee_I935 (.Y(N677), .A(a_man[22]), .B(b_man[22]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I960 (.Y(inst_cellmath__39[23]), .A(inst_cellmath__33[48]), .B(N4328));
XOR2XL inst_cellmath__45_0_I989 (.Y(N4562), .A(N677), .B(inst_cellmath__39[23]));
MX2XL cynw_cm_float_add2_ieee_I934 (.Y(N676), .A(a_man[21]), .B(b_man[21]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I959 (.Y(inst_cellmath__39[22]), .A(inst_cellmath__33[47]), .B(N4328));
XNOR2X1 inst_cellmath__45_0_I987 (.Y(N4508), .A(N676), .B(inst_cellmath__39[22]));
MX2XL cynw_cm_float_add2_ieee_I933 (.Y(N675), .A(a_man[20]), .B(b_man[20]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I958 (.Y(inst_cellmath__39[21]), .A(inst_cellmath__33[46]), .B(N4328));
XOR2XL inst_cellmath__45_0_I986 (.Y(N4581), .A(N675), .B(inst_cellmath__39[21]));
MX2XL cynw_cm_float_add2_ieee_I932 (.Y(N674), .A(a_man[19]), .B(b_man[19]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I957 (.Y(inst_cellmath__39[20]), .A(inst_cellmath__33[45]), .B(N4328));
XNOR2X1 inst_cellmath__45_0_I984 (.Y(N4521), .A(N674), .B(inst_cellmath__39[20]));
MX2XL cynw_cm_float_add2_ieee_I931 (.Y(N673), .A(a_man[18]), .B(b_man[18]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I956 (.Y(inst_cellmath__39[19]), .A(inst_cellmath__33[44]), .B(N4328));
XOR2XL inst_cellmath__45_0_I983 (.Y(N4599), .A(N673), .B(inst_cellmath__39[19]));
MX2XL cynw_cm_float_add2_ieee_I930 (.Y(N672), .A(a_man[17]), .B(b_man[17]), .S0(N3695));
XNOR2X1 inst_cellmath__39__19__2mx_I955 (.Y(inst_cellmath__39[18]), .A(inst_cellmath__33[43]), .B(N4328));
XNOR2X1 inst_cellmath__45_0_I981 (.Y(N4539), .A(N672), .B(inst_cellmath__39[18]));
NOR2XL inst_cellmath__45_0_I979 (.Y(N4588), .A(N671), .B(inst_cellmath__39[17]));
AOI21X4 inst_cellmath__45_0_I1006 (.Y(N4544), .A0(N4614), .A1(N4564), .B0(N4588));
OAI22X4 inst_cellmath__45_0_I1007 (.Y(N4512), .A0(N4539), .A1(N4544), .B0(inst_cellmath__39[18]), .B1(N672));
NOR2XL inst_cellmath__45_0_I982 (.Y(N4568), .A(N673), .B(inst_cellmath__39[19]));
AOI21X4 inst_cellmath__45_0_I1008 (.Y(N4605), .A0(N4599), .A1(N4512), .B0(N4568));
OAI22X4 inst_cellmath__45_0_I1009 (.Y(N4549), .A0(N4521), .A1(N4605), .B0(inst_cellmath__39[20]), .B1(N674));
NOR2XL inst_cellmath__45_0_I985 (.Y(N4550), .A(N675), .B(inst_cellmath__39[21]));
AOI21X4 inst_cellmath__45_0_I1010 (.Y(N4629), .A0(N4581), .A1(N4549), .B0(N4550));
OAI22X4 inst_cellmath__45_0_I1011 (.Y(N4558), .A0(N4508), .A1(N4629), .B0(inst_cellmath__39[22]), .B1(N676));
NOR2XL inst_cellmath__45_0_I988 (.Y(N4533), .A(N677), .B(inst_cellmath__39[23]));
AOI21X2 inst_cellmath__45_0_I1012 (.Y(N4622), .A0(N4562), .A1(N4558), .B0(N4533));
NOR2X1 inst_cellmath__45_0_I1038 (.Y(N4617), .A(inst_cellmath__39[24]), .B(N4622));
XOR2XL inst_cellmath__45_0_I2456 (.Y(N7112), .A(inst_cellmath__39[25]), .B(N4617));
CLKINVX1 inst_cellmath__62_0_I6953 (.Y(inst_cellmath__45[25]), .A(N7112));
XNOR2XL inst_cellmath__45_0_I1037 (.Y(inst_cellmath__45[24]), .A(inst_cellmath__39[24]), .B(N4622));
NOR2X2 inst_cellmath__49_0_I1071 (.Y(N4795), .A(inst_cellmath__45[24]), .B(inst_cellmath__45[25]));
XNOR2X1 inst_cellmath__45_0_I1036 (.Y(inst_cellmath__45[23]), .A(N4558), .B(N4562));
XNOR2X1 inst_cellmath__45_0_I1035 (.Y(inst_cellmath__45[22]), .A(N4629), .B(N4508));
NOR2X4 inst_cellmath__49_0_I1070 (.Y(N4773), .A(inst_cellmath__45[22]), .B(inst_cellmath__45[23]));
NAND2X4 inst_cellmath__49_0_I1084 (.Y(N4743), .A(N4773), .B(N4795));
XNOR2X1 inst_cellmath__45_0_I1034 (.Y(inst_cellmath__45[21]), .A(N4549), .B(N4581));
XNOR2X1 inst_cellmath__45_0_I1033 (.Y(inst_cellmath__45[20]), .A(N4605), .B(N4521));
NOR2XL inst_cellmath__49_0_I1066 (.Y(N4766), .A(inst_cellmath__45[21]), .B(inst_cellmath__45[20]));
XNOR2X1 inst_cellmath__45_0_I1032 (.Y(inst_cellmath__45[19]), .A(N4512), .B(N4599));
XNOR2X1 inst_cellmath__45_0_I1031 (.Y(inst_cellmath__45[18]), .A(N4544), .B(N4539));
NOR2XL inst_cellmath__49_0_I1065 (.Y(N4745), .A(inst_cellmath__45[19]), .B(inst_cellmath__45[18]));
NAND2X2 inst_cellmath__49_0_I1083 (.Y(N4724), .A(N4766), .B(N4745));
NOR2X4 inst_cellmath__49_0_I1091 (.Y(N4780), .A(N4724), .B(N4743));
NAND2X1 inst_cellmath__62_0_I6933 (.Y(N4729), .A(N4730), .B(N4780));
NAND2BXL inst_cellmath__49_0_I1075 (.Y(N4728), .AN(N4782), .B(N4802));
INVXL inst_cellmath__49_0_I1076 (.Y(N4747), .A(N4738));
AOI21XL inst_cellmath__49_0_I1077 (.Y(N4768), .A0(N4717), .A1(N4728), .B0(N4747));
NAND2BXL inst_cellmath__49_0_I1080 (.Y(N4756), .AN(N4745), .B(N4766));
INVXL inst_cellmath__49_0_I1081 (.Y(N4775), .A(N4795));
AOI21XL inst_cellmath__49_0_I1082 (.Y(N4797), .A0(N4773), .A1(N4756), .B0(N4775));
AOI21XL inst_cellmath__49_0_I1101 (.Y(N4750), .A0(N4780), .A1(N4768), .B0(N4797));
OAI21X1 cynw_cm_float_add2_ieee_I7125 (.Y(inst_cellmath__49[1]), .A0(N4784), .A1(N4729), .B0(N4750));
NAND2XL inst_cellmath__49_0_I1074 (.Y(N4779), .A(N4771), .B(N4752));
NAND2XL inst_cellmath__49_0_I1073 (.Y(N4760), .A(N4744), .B(N4725));
NAND2BXL inst_cellmath__49_0_I1085 (.Y(N4733), .AN(N4779), .B(N4760));
NOR2BX1 inst_cellmath__49_0_I1087 (.Y(N4761), .AN(N4788), .B(N4714));
INVXL inst_cellmath__49_0_I1088 (.Y(N4781), .A(N4743));
OAI21XL inst_cellmath__49_0_I1089 (.Y(N4801), .A0(N4724), .A1(N4761), .B0(N4781));
OA21X1 inst_cellmath__50_0_I2661 (.Y(N5079), .A0(N4729), .A1(N4733), .B0(N4801));
NOR2XL inst_cellmath__49_0_I1086 (.Y(N4719), .A(N4779), .B(N4760));
XOR2XL inst_cellmath__45_0_I1013 (.Y(inst_cellmath__45[0]), .A(inst_cellmath__44), .B(inst_cellmath__39[0]));
XNOR2X1 inst_cellmath__45_0_I1014 (.Y(inst_cellmath__45[1]), .A(N4556), .B(N4618));
NOR2BX1 inst_cellmath__49_0_I1040 (.Y(N4736), .AN(inst_cellmath__45[0]), .B(inst_cellmath__45[1]));
NOR2BX1 inst_cellmath__49_0_I1042 (.Y(N4757), .AN(inst_cellmath__45[2]), .B(inst_cellmath__45[3]));
INVXL inst_cellmath__49_0_I1043 (.Y(N4776), .A(inst_cellmath__45[5]));
OAI21XL inst_cellmath__49_0_I1044 (.Y(N4798), .A0(inst_cellmath__45[4]), .A1(N4757), .B0(N4776));
NOR2BX1 inst_cellmath__49_0_I1047 (.Y(N4786), .AN(inst_cellmath__45[6]), .B(inst_cellmath__45[7]));
INVXL inst_cellmath__49_0_I1048 (.Y(N4806), .A(inst_cellmath__45[9]));
OAI21XL inst_cellmath__49_0_I1049 (.Y(N4734), .A0(inst_cellmath__45[8]), .A1(N4786), .B0(N4806));
OAI21XL inst_cellmath__49_0_I1103 (.Y(N4723), .A0(N4779), .A1(N4798), .B0(N4734));
AOI21XL inst_cellmath__49_0_I1106 (.Y(N4751), .A0(N4719), .A1(N4736), .B0(N4723));
NOR2BX1 inst_cellmath__49_0_I1052 (.Y(N4720), .AN(inst_cellmath__45[10]), .B(inst_cellmath__45[11]));
INVXL inst_cellmath__49_0_I1053 (.Y(N4740), .A(inst_cellmath__45[13]));
OAI21XL inst_cellmath__49_0_I1054 (.Y(N4762), .A0(inst_cellmath__45[12]), .A1(N4720), .B0(N4740));
NOR2BX1 inst_cellmath__49_0_I1057 (.Y(N4748), .AN(inst_cellmath__45[14]), .B(inst_cellmath__45[15]));
INVXL inst_cellmath__49_0_I1058 (.Y(N4769), .A(inst_cellmath__45[17]));
OAI21XL inst_cellmath__49_0_I1059 (.Y(N4790), .A0(inst_cellmath__45[16]), .A1(N4748), .B0(N4769));
OAI21XL inst_cellmath__49_0_I1104 (.Y(N4765), .A0(N4714), .A1(N4762), .B0(N4790));
NOR2BX1 inst_cellmath__49_0_I1062 (.Y(N4777), .AN(inst_cellmath__45[18]), .B(inst_cellmath__45[19]));
INVXL inst_cellmath__49_0_I1063 (.Y(N4799), .A(inst_cellmath__45[21]));
OAI21XL inst_cellmath__49_0_I1064 (.Y(N4726), .A0(inst_cellmath__45[20]), .A1(N4777), .B0(N4799));
NOR2BX1 inst_cellmath__49_0_I1067 (.Y(N4712), .AN(inst_cellmath__45[22]), .B(inst_cellmath__45[23]));
INVXL inst_cellmath__49_0_I1068 (.Y(N4735), .A(inst_cellmath__45[25]));
OAI21XL inst_cellmath__49_0_I1069 (.Y(N4754), .A0(inst_cellmath__45[24]), .A1(N4712), .B0(N4735));
OAI21XL inst_cellmath__49_0_I1105 (.Y(N4805), .A0(N4726), .A1(N4743), .B0(N4754));
AOI21XL inst_cellmath__49_0_I1107 (.Y(N4793), .A0(N4780), .A1(N4765), .B0(N4805));
OA21X1 inst_cellmath__50_0_I2490 (.Y(N5135), .A0(N4751), .A1(N4729), .B0(N4793));
INVX2 inst_cellmath__50_0_I1198 (.Y(N5171), .A(N5135));
NOR2XL inst_cellmath__49_0_I1041 (.Y(N4715), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[0]));
NAND2BXL inst_cellmath__49_0_I1092 (.Y(N4789), .AN(N4715), .B(N4719));
INVX2 inst_cellmath__49_0_I1093 (.Y(N4716), .A(N4780));
AO21X4 inst_cellmath__50_0_I2658 (.Y(N5158), .A0(N4789), .A1(N4730), .B0(N4716));
AND2XL inst_cellmath__50_0_I1145 (.Y(N5031), .A(inst_cellmath__45[0]), .B(N5158));
NAND2XL inst_cellmath__62_0_I6932 (.Y(N4758), .A(N4715), .B(N4719));
NOR2BXL inst_cellmath__49_0_I1097 (.Y(inst_cellmath__49[4]), .AN(N4758), .B(N4729));
INVX8 inst_cellmath__50_0_I1170 (.Y(N5030), .A(inst_cellmath__49[4]));
NAND2X1 inst_cellmath__50_0_I1172 (.Y(N5022), .A(N5031), .B(N5030));
NOR2X2 inst_cellmath__50_0_I1199 (.Y(N5138), .A(N5022), .B(N5171));
NAND2X4 cynw_cm_float_add2_ieee_I7126 (.Y(N12575), .A(N5079), .B(N5138));
INVX3 inst_cellmath__50_0_I2594 (.Y(N7129), .A(N5158));
INVX2 inst_cellmath__50_0_I2600 (.Y(N7135), .A(N7129));
AND2XL inst_cellmath__50_0_I1147 (.Y(N5173), .A(inst_cellmath__45[2]), .B(N7135));
NAND2X1 inst_cellmath__50_0_I1174 (.Y(N5166), .A(N5173), .B(N5030));
AND2XL inst_cellmath__50_0_I1146 (.Y(N5102), .A(inst_cellmath__45[1]), .B(N7135));
NAND2XL inst_cellmath__50_0_I1173 (.Y(N5096), .A(N5030), .B(N5102));
AOI22X1 inst_cellmath__50_0_I1201 (.Y(N5117), .A0(N5135), .A1(N5166), .B0(N5171), .B1(N5096));
NAND2X2 cynw_cm_float_add2_ieee_I7127 (.Y(N5169), .A(N5079), .B(N5117));
INVX3 cynw_cm_float_add2_ieee_I7128 (.Y(N5023), .A(inst_cellmath__49[1]));
INVX2 cynw_cm_float_add2_ieee_I7129 (.Y(N5059), .A(N5023));
AOI22X2 cynw_cm_float_add2_ieee_I7130 (.Y(inst_cellmath__50[2]), .A0(N5059), .A1(N12575), .B0(N5023), .B1(N5169));
NAND2XL hyperpropagate_3_1_A_I7335 (.Y(N12741), .A(N12585), .B(rm[0]));
NOR2XL hyperpropagate_3_1_A_I7336 (.Y(inst_cellmath__5), .A(rm[1]), .B(N12741));
INVXL cynw_cm_float_add2_ieee_I7133 (.Y(N5354), .A(inst_cellmath__48));
AND2XL cynw_cm_float_add2_ieee_I7134 (.Y(N635), .A(inst_cellmath__5), .B(N5354));
AND2XL cynw_cm_float_add2_ieee_I7135 (.Y(N634), .A(inst_cellmath__6), .B(inst_cellmath__48));
NOR3BXL cynw_cm_float_add2_ieee_I7136 (.Y(inst_cellmath__8), .AN(N12547), .B(N12585), .C(rm[0]));
NOR3XL cynw_cm_float_add2_ieee_I7137 (.Y(inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
INVXL cynw_cm_float_add2_ieee_I7138 (.Y(N12558), .A(inst_cellmath__49[1]));
OR2XL cynw_cm_float_add2_ieee_I1281 (.Y(N628), .A(inst_cellmath__33[24]), .B(inst_cellmath__42));
XNOR2X1 cynw_cm_float_add2_ieee_I1278 (.Y(N626), .A(inst_cellmath__42), .B(inst_cellmath__33[24]));
OR2XL cynw_cm_float_add2_ieee_I1280 (.Y(N627), .A(inst_cellmath__30), .B(N626));
OAI2BB1X1 cynw_cm_float_add2_ieee_I2663 (.Y(N630), .A0N(inst_cellmath__30), .A1N(N628), .B0(N627));
MX2XL cynw_cm_float_add2_ieee_I1284 (.Y(inst_cellmath__43), .A(inst_cellmath__33[24]), .B(N630), .S0(inst_cellmath__39[25]));
NOR2XL cynw_cm_float_add2_ieee_I1292 (.Y(N5374), .A(inst_cellmath__42), .B(inst_cellmath__43));
OAI21X2 cynw_cm_float_add2_ieee_I7140 (.Y(N12567), .A0(N5059), .A1(N12575), .B0(N5374));
MX2XL cynw_cm_float_add2_ieee_I7141 (.Y(inst_cellmath__54), .A(inst_cellmath__42), .B(N12567), .S0(N12558));
OAI21XL cynw_cm_float_add2_ieee_I7142 (.Y(N12573), .A0(N12548), .A1(N12565), .B0(inst_cellmath__6));
NOR2BX1 cynw_cm_float_add2_ieee_I7143 (.Y(N12557), .AN(N12573), .B(inst_cellmath__8));
INVX2 cynw_cm_float_add2_ieee_I7144 (.Y(N12592), .A(inst_cellmath__50[2]));
MXI2X1 cynw_cm_float_add2_ieee_I7145 (.Y(N12550), .A(inst_cellmath__42), .B(N12567), .S0(N12558));
NAND2X2 cynw_cm_float_add2_ieee_I7146 (.Y(N12560), .A(N12550), .B(N12592));
AOI21X2 cynw_cm_float_add2_ieee_I7147 (.Y(N12578), .A0(inst_cellmath__4), .A1(N12560), .B0(N635));
NAND2X1 cynw_cm_float_add2_ieee_I7148 (.Y(N636), .A(N12557), .B(N12578));
NOR2XL inst_cellmath__62_0_I6934 (.Y(inst_cellmath__49[5]), .A(N4758), .B(N4729));
OR2XL cmp_A_I7337 (.Y(N12748), .A(a_sign), .B(b_sign));
AO22XL cmp_A_I7338 (.Y(N645), .A0(N12748), .A1(inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL cynw_cm_float_add2_ieee_I1114 (.Y(inst_cellmath__66), .A(inst_cellmath__11), .B(inst_cellmath__16), .C(N645));
NOR2BX1 inst_cellmath__64__48__2WWMM_I1115 (.Y(N4931), .AN(inst_cellmath__18), .B(inst_cellmath__13));
AOI22XL inst_cellmath__64__48__2WWMM_I1116 (.Y(N4952), .A0(a_sign), .A1(inst_cellmath__13), .B0(N4931), .B1(b_sign));
AO22XL inst_cellmath__64__48__2WWMM_I1117 (.Y(inst_cellmath__64[0]), .A0(inst_cellmath__13), .A1(N11653), .B0(N4931), .B1(b_man[0]));
AO22XL inst_cellmath__64__48__2WWMM_I1118 (.Y(inst_cellmath__64[1]), .A0(inst_cellmath__13), .A1(a_man[1]), .B0(N4931), .B1(b_man[1]));
AO22XL inst_cellmath__64__48__2WWMM_I1119 (.Y(inst_cellmath__64[2]), .A0(inst_cellmath__13), .A1(a_man[2]), .B0(N4931), .B1(b_man[2]));
AO22XL inst_cellmath__64__48__2WWMM_I1120 (.Y(inst_cellmath__64[3]), .A0(inst_cellmath__13), .A1(a_man[3]), .B0(N4931), .B1(b_man[3]));
AO22XL inst_cellmath__64__48__2WWMM_I1121 (.Y(inst_cellmath__64[4]), .A0(inst_cellmath__13), .A1(a_man[4]), .B0(N4931), .B1(b_man[4]));
AO22XL inst_cellmath__64__48__2WWMM_I1122 (.Y(inst_cellmath__64[5]), .A0(inst_cellmath__13), .A1(a_man[5]), .B0(N4931), .B1(b_man[5]));
AO22XL inst_cellmath__64__48__2WWMM_I1123 (.Y(inst_cellmath__64[6]), .A0(inst_cellmath__13), .A1(a_man[6]), .B0(N4931), .B1(b_man[6]));
AO22XL inst_cellmath__64__48__2WWMM_I1124 (.Y(inst_cellmath__64[7]), .A0(inst_cellmath__13), .A1(a_man[7]), .B0(N4931), .B1(b_man[7]));
AO22XL inst_cellmath__64__48__2WWMM_I1125 (.Y(inst_cellmath__64[8]), .A0(inst_cellmath__13), .A1(a_man[8]), .B0(N4931), .B1(b_man[8]));
AO22XL inst_cellmath__64__48__2WWMM_I1126 (.Y(inst_cellmath__64[9]), .A0(inst_cellmath__13), .A1(a_man[9]), .B0(N4931), .B1(b_man[9]));
AO22XL inst_cellmath__64__48__2WWMM_I1127 (.Y(inst_cellmath__64[10]), .A0(inst_cellmath__13), .A1(a_man[10]), .B0(N4931), .B1(b_man[10]));
AO22XL inst_cellmath__64__48__2WWMM_I1128 (.Y(inst_cellmath__64[11]), .A0(inst_cellmath__13), .A1(a_man[11]), .B0(N4931), .B1(b_man[11]));
AO22XL inst_cellmath__64__48__2WWMM_I1129 (.Y(inst_cellmath__64[12]), .A0(inst_cellmath__13), .A1(a_man[12]), .B0(N4931), .B1(b_man[12]));
AO22XL inst_cellmath__64__48__2WWMM_I1130 (.Y(inst_cellmath__64[13]), .A0(inst_cellmath__13), .A1(a_man[13]), .B0(N4931), .B1(b_man[13]));
AO22XL inst_cellmath__64__48__2WWMM_I1131 (.Y(inst_cellmath__64[14]), .A0(inst_cellmath__13), .A1(a_man[14]), .B0(N4931), .B1(b_man[14]));
AO22XL inst_cellmath__64__48__2WWMM_I1132 (.Y(inst_cellmath__64[15]), .A0(inst_cellmath__13), .A1(a_man[15]), .B0(N4931), .B1(b_man[15]));
AO22XL inst_cellmath__64__48__2WWMM_I1133 (.Y(inst_cellmath__64[16]), .A0(inst_cellmath__13), .A1(a_man[16]), .B0(N4931), .B1(b_man[16]));
AO22XL inst_cellmath__64__48__2WWMM_I1134 (.Y(inst_cellmath__64[17]), .A0(inst_cellmath__13), .A1(a_man[17]), .B0(N4931), .B1(b_man[17]));
AO22XL inst_cellmath__64__48__2WWMM_I1135 (.Y(inst_cellmath__64[18]), .A0(inst_cellmath__13), .A1(a_man[18]), .B0(N4931), .B1(b_man[18]));
AO22XL inst_cellmath__64__48__2WWMM_I1136 (.Y(inst_cellmath__64[19]), .A0(inst_cellmath__13), .A1(a_man[19]), .B0(N4931), .B1(b_man[19]));
AO22XL inst_cellmath__64__48__2WWMM_I1137 (.Y(inst_cellmath__64[20]), .A0(inst_cellmath__13), .A1(a_man[20]), .B0(N4931), .B1(b_man[20]));
AO22XL inst_cellmath__64__48__2WWMM_I1138 (.Y(inst_cellmath__64[21]), .A0(inst_cellmath__13), .A1(a_man[21]), .B0(N4931), .B1(b_man[21]));
OAI21XL inst_cellmath__64__48__2WWMM_I1139 (.Y(N710), .A0(inst_cellmath__18), .A1(inst_cellmath__13), .B0(N4952));
OR3X1 inst_cellmath__62_0_I6930 (.Y(inst_cellmath__63), .A(inst_cellmath__13), .B(inst_cellmath__18), .C(N547));
MX2XL inst_cellmath__67_0_I1140 (.Y(N5001), .A(inst_cellmath__66), .B(N710), .S0(inst_cellmath__63));
AND2XL inst_cellmath__62_0_I6931 (.Y(N706), .A(inst_cellmath__11), .B(inst_cellmath__16));
NOR2XL inst_cellmath__67_0_I1141 (.Y(N5010), .A(inst_cellmath__63), .B(N706));
MX2XL inst_cellmath__67_0_I7231 (.Y(N5004), .A(inst_cellmath__48), .B(inst_cellmath__6), .S0(inst_cellmath__49[5]));
MX2XL inst_cellmath__67_0_I1143 (.Y(x[31]), .A(N5001), .B(N5004), .S0(N5010));
INVXL inst_cellmath__50_0_I2599 (.Y(N7134), .A(N7129));
AND2XL inst_cellmath__50_0_I1148 (.Y(N5080), .A(N7135), .B(inst_cellmath__45[3]));
AND2XL inst_cellmath__50_0_I1149 (.Y(N5151), .A(N7135), .B(inst_cellmath__45[4]));
AND2XL inst_cellmath__50_0_I1150 (.Y(N5060), .A(N7134), .B(inst_cellmath__45[5]));
AND2XL inst_cellmath__50_0_I1151 (.Y(N5130), .A(N7134), .B(inst_cellmath__45[6]));
AND2XL inst_cellmath__50_0_I1152 (.Y(N5040), .A(N7134), .B(inst_cellmath__45[7]));
MX2XL inst_cellmath__50_0_I1153 (.Y(N5111), .A(inst_cellmath__45[0]), .B(inst_cellmath__45[8]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1154 (.Y(N5146), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[9]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1155 (.Y(N5016), .A(inst_cellmath__45[2]), .B(inst_cellmath__45[10]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1156 (.Y(N5053), .A(inst_cellmath__45[3]), .B(inst_cellmath__45[11]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1157 (.Y(N5090), .A(inst_cellmath__45[4]), .B(inst_cellmath__45[12]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1158 (.Y(N5124), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[13]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1159 (.Y(N5160), .A(inst_cellmath__45[6]), .B(inst_cellmath__45[14]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1160 (.Y(N5034), .A(inst_cellmath__45[7]), .B(inst_cellmath__45[15]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1161 (.Y(N5068), .A(inst_cellmath__45[8]), .B(inst_cellmath__45[16]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1162 (.Y(N5105), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[17]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1163 (.Y(N5139), .A(inst_cellmath__45[10]), .B(inst_cellmath__45[18]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1164 (.Y(N5176), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[19]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1165 (.Y(N5047), .A(inst_cellmath__45[12]), .B(inst_cellmath__45[20]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1166 (.Y(N5084), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[21]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1167 (.Y(N5119), .A(inst_cellmath__45[14]), .B(inst_cellmath__45[22]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1168 (.Y(N5155), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[23]), .S0(N7134));
MX2XL inst_cellmath__50_0_I1169 (.Y(N5026), .A(inst_cellmath__45[16]), .B(inst_cellmath__45[24]), .S0(N7134));
INVXL inst_cellmath__50_0_I1171 (.Y(N5066), .A(N5030));
NAND2XL inst_cellmath__50_0_I1175 (.Y(N5074), .A(N5080), .B(N5030));
NAND2XL inst_cellmath__50_0_I1176 (.Y(N5145), .A(N5151), .B(N5030));
NAND2XL inst_cellmath__50_0_I1177 (.Y(N5052), .A(N5060), .B(N5030));
NAND2XL inst_cellmath__50_0_I1178 (.Y(N5123), .A(N5130), .B(N5030));
NAND2XL inst_cellmath__50_0_I1179 (.Y(N5033), .A(N5040), .B(N5030));
NAND2XL inst_cellmath__50_0_I1180 (.Y(N5104), .A(N5111), .B(N5030));
NAND2XL inst_cellmath__50_0_I1181 (.Y(N5175), .A(N5146), .B(N5030));
NAND2XL inst_cellmath__50_0_I1182 (.Y(N5083), .A(N5016), .B(N5030));
NAND2XL inst_cellmath__50_0_I1183 (.Y(N5154), .A(N5053), .B(N5030));
NAND2XL inst_cellmath__50_0_I1184 (.Y(N5063), .A(N5090), .B(N5030));
NAND2XL inst_cellmath__50_0_I1185 (.Y(N5133), .A(N5124), .B(N5030));
NAND2XL inst_cellmath__50_0_I1186 (.Y(N5043), .A(N5160), .B(N5030));
NAND2XL inst_cellmath__50_0_I1187 (.Y(N5114), .A(N5034), .B(N5030));
AOI22XL inst_cellmath__50_0_I1188 (.Y(N5019), .A0(N5031), .A1(N5066), .B0(N5068), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1189 (.Y(N5056), .A0(N5102), .A1(N5066), .B0(N5105), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1190 (.Y(N5093), .A0(N5173), .A1(N5066), .B0(N5139), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1191 (.Y(N5127), .A0(N5080), .A1(N5066), .B0(N5176), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1192 (.Y(N5163), .A0(N5151), .A1(N5066), .B0(N5047), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1193 (.Y(N5037), .A0(N5066), .A1(N5060), .B0(N5084), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1194 (.Y(N5071), .A0(N5066), .A1(N5130), .B0(N5119), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1195 (.Y(N5108), .A0(N5066), .A1(N5040), .B0(N5155), .B1(N5030));
AOI22XL inst_cellmath__50_0_I1196 (.Y(N5142), .A0(N5066), .A1(N5111), .B0(N5026), .B1(N5030));
INVXL inst_cellmath__50_0_I6631 (.Y(N11648), .A(N5135));
INVX1 inst_cellmath__50_0_I6632 (.Y(N11649), .A(N11648));
INVXL inst_cellmath__50_0_I6731 (.Y(N11788), .A(N11649));
INVX1 inst_cellmath__50_0_I6732 (.Y(N11789), .A(N11788));
INVX1 inst_cellmath__50_0_I6633 (.Y(N11650), .A(N5171));
INVX3 inst_cellmath__50_0_I6634 (.Y(N11651), .A(N11650));
AOI22XL inst_cellmath__50_0_I1200 (.Y(N5081), .A0(N5096), .A1(N11649), .B0(N11651), .B1(N5022));
AOI22XL inst_cellmath__50_0_I1202 (.Y(N5153), .A0(N5074), .A1(N11789), .B0(N5166), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1203 (.Y(N5025), .A0(N11789), .A1(N5145), .B0(N5074), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1204 (.Y(N5062), .A0(N11789), .A1(N5052), .B0(N5145), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1205 (.Y(N5098), .A0(N11789), .A1(N5123), .B0(N5052), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1206 (.Y(N5131), .A0(N11789), .A1(N5033), .B0(N5123), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1207 (.Y(N5167), .A0(N11789), .A1(N5104), .B0(N5033), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1208 (.Y(N5042), .A0(N11789), .A1(N5175), .B0(N5104), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1209 (.Y(N5076), .A0(N11789), .A1(N5083), .B0(N5175), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1210 (.Y(N5113), .A0(N11789), .A1(N5154), .B0(N5083), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1211 (.Y(N5148), .A0(N11789), .A1(N5063), .B0(N5154), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1212 (.Y(N5017), .A0(N11789), .A1(N5133), .B0(N5063), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1213 (.Y(N5054), .A0(N11789), .A1(N5043), .B0(N5133), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1214 (.Y(N5092), .A0(N11789), .A1(N5114), .B0(N5043), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1215 (.Y(N5126), .A0(N11789), .A1(N5019), .B0(N5114), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1216 (.Y(N5162), .A0(N11789), .A1(N5056), .B0(N5019), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1217 (.Y(N5036), .A0(N11789), .A1(N5093), .B0(N5056), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1218 (.Y(N5069), .A0(N11789), .A1(N5127), .B0(N5093), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1219 (.Y(N5106), .A0(N11789), .A1(N5163), .B0(N5127), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1220 (.Y(N5141), .A0(N11789), .A1(N5037), .B0(N5163), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1221 (.Y(N5178), .A0(N11789), .A1(N5071), .B0(N5037), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1222 (.Y(N5049), .A0(N11789), .A1(N5108), .B0(N5071), .B1(N11651));
AOI22XL inst_cellmath__50_0_I1223 (.Y(N5086), .A0(N11789), .A1(N5142), .B0(N5108), .B1(N11651));
INVXL inst_cellmath__50_0_I1225 (.Y(N5116), .A(N5079));
NAND2X1 inst_cellmath__50_0_I1227 (.Y(N5099), .A(N5079), .B(N5081));
NAND2XL inst_cellmath__50_0_I1229 (.Y(N5077), .A(N5153), .B(N5079));
AOI22XL inst_cellmath__50_0_I1230 (.Y(N5149), .A0(N5116), .A1(N5138), .B0(N5025), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1231 (.Y(N5020), .A0(N5116), .A1(N5081), .B0(N5062), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1232 (.Y(N5057), .A0(N5116), .A1(N5117), .B0(N5098), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1233 (.Y(N5094), .A0(N5116), .A1(N5153), .B0(N5131), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1234 (.Y(N5128), .A0(N5116), .A1(N5025), .B0(N5167), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1235 (.Y(N5164), .A0(N5116), .A1(N5062), .B0(N5042), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1236 (.Y(N5038), .A0(N5116), .A1(N5098), .B0(N5076), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1237 (.Y(N5072), .A0(N5116), .A1(N5131), .B0(N5113), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1238 (.Y(N5109), .A0(N5116), .A1(N5167), .B0(N5148), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1239 (.Y(N5143), .A0(N5116), .A1(N5042), .B0(N5017), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1240 (.Y(N5179), .A0(N5116), .A1(N5076), .B0(N5054), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1241 (.Y(N5050), .A0(N5116), .A1(N5113), .B0(N5092), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1242 (.Y(N5087), .A0(N5116), .A1(N5148), .B0(N5126), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1243 (.Y(N5121), .A0(N5116), .A1(N5017), .B0(N5162), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1244 (.Y(N5157), .A0(N5116), .A1(N5054), .B0(N5036), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1245 (.Y(N5029), .A0(N5116), .A1(N5092), .B0(N5069), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1246 (.Y(N5065), .A0(N5116), .A1(N5126), .B0(N5106), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1247 (.Y(N5101), .A0(N5116), .A1(N5162), .B0(N5141), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1248 (.Y(N5136), .A0(N5116), .A1(N5036), .B0(N5178), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1249 (.Y(N5172), .A0(N5116), .A1(N5069), .B0(N5049), .B1(N5079));
AOI22XL inst_cellmath__50_0_I1250 (.Y(N5045), .A0(N5116), .A1(N5106), .B0(N5086), .B1(N5079));
NOR2XL inst_cellmath__50_0_I1254 (.Y(inst_cellmath__50[1]), .A(N5059), .B(N5099));
AOI22XL inst_cellmath__50_0_I1256 (.Y(inst_cellmath__50[3]), .A0(N5023), .A1(N5077), .B0(N5099), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1257 (.Y(inst_cellmath__50[4]), .A0(N5023), .A1(N5149), .B0(N5169), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1258 (.Y(inst_cellmath__50[5]), .A0(N5023), .A1(N5020), .B0(N5077), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1259 (.Y(inst_cellmath__50[6]), .A0(N5023), .A1(N5057), .B0(N5149), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1260 (.Y(inst_cellmath__50[7]), .A0(N5023), .A1(N5094), .B0(N5020), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1261 (.Y(inst_cellmath__50[8]), .A0(N5023), .A1(N5128), .B0(N5057), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1262 (.Y(inst_cellmath__50[9]), .A0(N5023), .A1(N5164), .B0(N5094), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1263 (.Y(inst_cellmath__50[10]), .A0(N5023), .A1(N5038), .B0(N5128), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1264 (.Y(inst_cellmath__50[11]), .A0(N5023), .A1(N5072), .B0(N5164), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1265 (.Y(inst_cellmath__50[12]), .A0(N5023), .A1(N5109), .B0(N5038), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1266 (.Y(inst_cellmath__50[13]), .A0(N5023), .A1(N5143), .B0(N5072), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1267 (.Y(inst_cellmath__50[14]), .A0(N5023), .A1(N5179), .B0(N5109), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1268 (.Y(inst_cellmath__50[15]), .A0(N5023), .A1(N5050), .B0(N5143), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1269 (.Y(inst_cellmath__50[16]), .A0(N5023), .A1(N5087), .B0(N5179), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1270 (.Y(inst_cellmath__50[17]), .A0(N5023), .A1(N5121), .B0(N5050), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1271 (.Y(inst_cellmath__50[18]), .A0(N5023), .A1(N5157), .B0(N5087), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1272 (.Y(inst_cellmath__50[19]), .A0(N5023), .A1(N5029), .B0(N5121), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1273 (.Y(inst_cellmath__50[20]), .A0(N5023), .A1(N5065), .B0(N5157), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1274 (.Y(inst_cellmath__50[21]), .A0(N5023), .A1(N5101), .B0(N5029), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1275 (.Y(inst_cellmath__50[22]), .A0(N5023), .A1(N5136), .B0(N5065), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1276 (.Y(inst_cellmath__50[23]), .A0(N5023), .A1(N5172), .B0(N5101), .B1(N5059));
AOI22XL inst_cellmath__50_0_I1277 (.Y(inst_cellmath__50[24]), .A0(N5023), .A1(N5045), .B0(N5136), .B1(N5059));
MX2XL cynw_cm_float_add2_ieee_I1285 (.Y(inst_cellmath__53), .A(inst_cellmath__50[1]), .B(inst_cellmath__43), .S0(inst_cellmath__49[1]));
OAI21X2 cynw_cm_float_add2_ieee_I2709 (.Y(N639), .A0(N634), .A1(N635), .B0(inst_cellmath__54));
OAI2BB1XL cynw_cm_float_add2_ieee_I2494 (.Y(inst_cellmath__55), .A0N(inst_cellmath__53), .A1N(N636), .B0(N639));
ADDHXL inst_cellmath__57_0_I1302 (.CO(N5477), .S(inst_cellmath__57[0]), .A(inst_cellmath__50[2]), .B(inst_cellmath__55));
ADDHXL inst_cellmath__57_0_I1303 (.CO(N5466), .S(inst_cellmath__57[1]), .A(inst_cellmath__50[3]), .B(N5477));
ADDHXL inst_cellmath__57_0_I1304 (.CO(N5456), .S(inst_cellmath__57[2]), .A(inst_cellmath__50[4]), .B(N5466));
ADDHXL inst_cellmath__57_0_I1305 (.CO(N5449), .S(inst_cellmath__57[3]), .A(inst_cellmath__50[5]), .B(N5456));
ADDHXL inst_cellmath__57_0_I1306 (.CO(N5438), .S(inst_cellmath__57[4]), .A(inst_cellmath__50[6]), .B(N5449));
ADDHXL inst_cellmath__57_0_I1307 (.CO(N5429), .S(inst_cellmath__57[5]), .A(inst_cellmath__50[7]), .B(N5438));
ADDHXL inst_cellmath__57_0_I1308 (.CO(N5421), .S(inst_cellmath__57[6]), .A(inst_cellmath__50[8]), .B(N5429));
ADDHXL inst_cellmath__57_0_I1309 (.CO(N5482), .S(inst_cellmath__57[7]), .A(inst_cellmath__50[9]), .B(N5421));
ADDHXL inst_cellmath__57_0_I1310 (.CO(N5474), .S(inst_cellmath__57[8]), .A(inst_cellmath__50[10]), .B(N5482));
ADDHXL inst_cellmath__57_0_I1311 (.CO(N5464), .S(inst_cellmath__57[9]), .A(inst_cellmath__50[11]), .B(N5474));
ADDHXL inst_cellmath__57_0_I1312 (.CO(N5454), .S(inst_cellmath__57[10]), .A(inst_cellmath__50[12]), .B(N5464));
ADDHXL inst_cellmath__57_0_I1313 (.CO(N5446), .S(inst_cellmath__57[11]), .A(inst_cellmath__50[13]), .B(N5454));
ADDHXL inst_cellmath__57_0_I1314 (.CO(N5436), .S(inst_cellmath__57[12]), .A(inst_cellmath__50[14]), .B(N5446));
ADDHXL inst_cellmath__57_0_I1315 (.CO(N5428), .S(inst_cellmath__57[13]), .A(inst_cellmath__50[15]), .B(N5436));
ADDHXL inst_cellmath__57_0_I1316 (.CO(N5418), .S(inst_cellmath__57[14]), .A(inst_cellmath__50[16]), .B(N5428));
ADDHXL inst_cellmath__57_0_I1317 (.CO(N5480), .S(inst_cellmath__57[15]), .A(inst_cellmath__50[17]), .B(N5418));
ADDHXL inst_cellmath__57_0_I1318 (.CO(N5473), .S(inst_cellmath__57[16]), .A(inst_cellmath__50[18]), .B(N5480));
ADDHXL inst_cellmath__57_0_I1319 (.CO(N5461), .S(inst_cellmath__57[17]), .A(inst_cellmath__50[19]), .B(N5473));
ADDHXL inst_cellmath__57_0_I1320 (.CO(N5452), .S(inst_cellmath__57[18]), .A(inst_cellmath__50[20]), .B(N5461));
ADDHXL inst_cellmath__57_0_I1321 (.CO(N5445), .S(inst_cellmath__57[19]), .A(inst_cellmath__50[21]), .B(N5452));
ADDHXL inst_cellmath__57_0_I1322 (.CO(N5434), .S(inst_cellmath__57[20]), .A(inst_cellmath__50[22]), .B(N5445));
ADDHXL inst_cellmath__57_0_I1323 (.CO(N5426), .S(inst_cellmath__57[21]), .A(inst_cellmath__50[23]), .B(N5434));
ADDHXL inst_cellmath__57_0_I1324 (.CO(inst_cellmath__57[23]), .S(inst_cellmath__57[22]), .A(inst_cellmath__50[24]), .B(N5426));
INVXL cynw_cm_float_add2_ieee_I76 (.Y(N574), .A(N3367));
MX2XL inst_cellmath__29_0_I1327 (.Y(inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(N574));
MX2XL inst_cellmath__29_0_I1328 (.Y(inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(N574));
MX2XL inst_cellmath__29_0_I1329 (.Y(inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(N574));
MX2XL inst_cellmath__29_0_I1330 (.Y(inst_cellmath__29[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(N574));
MX2XL inst_cellmath__29_0_I1331 (.Y(inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(N574));
MX2XL inst_cellmath__29_0_I1332 (.Y(inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(N574));
MX2XL inst_cellmath__29_0_I1333 (.Y(inst_cellmath__29[6]), .A(a_exp[6]), .B(b_exp[6]), .S0(N574));
MX2XL inst_cellmath__62_0_I6936 (.Y(inst_cellmath__29[7]), .A(a_exp[7]), .B(b_exp[7]), .S0(N574));
NAND3XL inst_cellmath__62_0_I1336 (.Y(N5584), .A(inst_cellmath__29[6]), .B(inst_cellmath__29[7]), .C(inst_cellmath__29[5]));
NOR2XL inst_cellmath__62_0_I1337 (.Y(N5583), .A(inst_cellmath__29[0]), .B(N5584));
NAND3XL inst_cellmath__62_0_I1338 (.Y(N5580), .A(inst_cellmath__29[4]), .B(inst_cellmath__29[3]), .C(N5583));
AND2XL inst_cellmath__62_0_I6935 (.Y(N12151), .A(inst_cellmath__45[24]), .B(inst_cellmath__57[23]));
ADDFXL inst_cellmath__62_0_I6937 (.CO(N12123), .S(inst_cellmath__59[0]), .A(N5135), .B(inst_cellmath__29[0]), .CI(inst_cellmath__57[23]));
INVXL cynw_cm_float_add2_ieee_I1346 (.Y(N5614), .A(inst_cellmath__29[1]));
ADDFHXL inst_cellmath__62_0_I6938 (.CO(N12160), .S(inst_cellmath__59[1]), .A(N5614), .B(N5023), .CI(N12123));
ADDHX1 cynw_cm_float_add2_ieee_I1347 (.CO(N5619), .S(N5605), .A(inst_cellmath__29[1]), .B(inst_cellmath__29[2]));
ADDFHXL inst_cellmath__62_0_I6939 (.CO(N12194), .S(inst_cellmath__59[2]), .A(N5079), .B(N5605), .CI(N12160));
ADDHX1 cynw_cm_float_add2_ieee_I1348 (.CO(N5592), .S(N5630), .A(inst_cellmath__29[3]), .B(N5619));
ADDFHXL inst_cellmath__62_0_I6940 (.CO(N12148), .S(inst_cellmath__59[3]), .A(N5158), .B(N5630), .CI(N12194));
ADDHX1 cynw_cm_float_add2_ieee_I1349 (.CO(N5612), .S(N5600), .A(inst_cellmath__29[4]), .B(N5592));
ADDFHXL inst_cellmath__62_0_I6941 (.CO(N12184), .S(inst_cellmath__59[4]), .A(N5030), .B(N5600), .CI(N12148));
INVXL cynw_cm_float_add2_ieee_I1350 (.Y(N5622), .A(inst_cellmath__29[5]));
ADDFHXL inst_cellmath__62_0_I6942 (.CO(N12139), .S(inst_cellmath__59[5]), .A(N5612), .B(N5622), .CI(N12184));
INVXL cynw_cm_float_add2_ieee_I1351 (.Y(N5617), .A(inst_cellmath__29[6]));
ADDFHXL inst_cellmath__62_0_I6943 (.CO(N12174), .S(inst_cellmath__59[6]), .A(N5617), .B(inst_cellmath__29[5]), .CI(N12139));
INVXL cynw_cm_float_add2_ieee_I1352 (.Y(N5610), .A(inst_cellmath__29[7]));
ADDFHXL inst_cellmath__62_0_I6944 (.CO(N12129), .S(inst_cellmath__59[7]), .A(N5610), .B(inst_cellmath__29[6]), .CI(N12174));
XNOR2X1 inst_cellmath__62_0_I6945 (.Y(N12145), .A(inst_cellmath__29[7]), .B(N12129));
NOR2XL inst_cellmath__62_0_I6946 (.Y(N12165), .A(inst_cellmath__29[7]), .B(N12129));
OR3XL inst_cellmath__62_0_I7276 (.Y(N12188), .A(inst_cellmath__59[0]), .B(inst_cellmath__59[1]), .C(inst_cellmath__59[3]));
NOR3X2 inst_cellmath__62_0_I6951 (.Y(N12177), .A(N12188), .B(inst_cellmath__59[7]), .C(N12145));
OR4X1 inst_cellmath__62_0_I6952 (.Y(N12189), .A(N706), .B(inst_cellmath__17), .C(inst_cellmath__12), .D(inst_cellmath__63));
NAND3BXL inst_cellmath__62_0_I6954 (.Y(N12134), .AN(N5580), .B(inst_cellmath__29[1]), .C(inst_cellmath__29[2]));
NOR2XL andori2bb1_A_I7339 (.Y(N12755), .A(N12151), .B(inst_cellmath__45[25]));
NOR2XL andori2bb1_A_I7340 (.Y(inst_cellmath__62), .A(N12755), .B(N12134));
NOR4X1 inst_cellmath__62_0_I6956 (.Y(N12125), .A(N12189), .B(inst_cellmath__49[5]), .C(inst_cellmath__62), .D(N12165));
NOR4X1 inst_cellmath__62_0_I7236 (.Y(N12157), .A(inst_cellmath__59[2]), .B(inst_cellmath__59[4]), .C(inst_cellmath__59[5]), .D(inst_cellmath__59[6]));
NAND2X1 inst_cellmath__62_0_I6959 (.Y(N12162), .A(N12157), .B(N12177));
NAND2X1 inst_cellmath__62_0_I6960 (.Y(inst_cellmath__71), .A(N12125), .B(N12162));
OR4X1 cynw_cm_float_add2_ieee_I2668 (.Y(N650), .A(inst_cellmath__4), .B(inst_cellmath__8), .C(N634), .D(N635));
AND2XL cynw_cm_float_add2_ieee_I1375 (.Y(N651), .A(N650), .B(inst_cellmath__62));
OR4X1 cynw_cm_float_add2_ieee_I1376 (.Y(inst_cellmath__68[0]), .A(inst_cellmath__17), .B(inst_cellmath__12), .C(inst_cellmath__63), .D(N651));
OR4X1 inst_cellmath__72_0_I2669 (.Y(N5745), .A(inst_cellmath__12), .B(inst_cellmath__17), .C(inst_cellmath__63), .D(inst_cellmath__62));
INVX3 inst_cellmath__72_0_I1380 (.Y(N5751), .A(inst_cellmath__71));
INVXL inst_cellmath__72_0_I1381 (.Y(N5733), .A(N5751));
MX2XL inst_cellmath__72_0_I1382 (.Y(x[23]), .A(inst_cellmath__59[0]), .B(inst_cellmath__68[0]), .S0(N5733));
MX2XL inst_cellmath__72_0_I1383 (.Y(x[24]), .A(inst_cellmath__59[1]), .B(N5745), .S0(N5733));
MX2XL inst_cellmath__72_0_I1384 (.Y(x[25]), .A(inst_cellmath__59[2]), .B(N5745), .S0(N5733));
MX2XL inst_cellmath__72_0_I1385 (.Y(x[26]), .A(inst_cellmath__59[3]), .B(N5745), .S0(N5733));
MX2XL inst_cellmath__72_0_I1386 (.Y(x[27]), .A(inst_cellmath__59[4]), .B(N5745), .S0(N5733));
MX2XL inst_cellmath__72_0_I1387 (.Y(x[28]), .A(inst_cellmath__59[5]), .B(N5745), .S0(N5733));
MX2XL inst_cellmath__72_0_I1388 (.Y(x[29]), .A(inst_cellmath__59[6]), .B(N5745), .S0(N5733));
MX2XL inst_cellmath__72_0_I1389 (.Y(x[30]), .A(inst_cellmath__59[7]), .B(N5745), .S0(N5733));
NAND2XL inst_cellmath__7_0_I1390 (.Y(N5769), .A(rm[0]), .B(rm[1]));
NOR2XL inst_cellmath__7_0_I1391 (.Y(inst_cellmath__7), .A(rm[2]), .B(N5769));
MXI2XL cynw_cm_float_add2_ieee_I1393 (.Y(N652), .A(inst_cellmath__48), .B(N5354), .S0(inst_cellmath__5));
OR2XL cynw_cm_float_add2_ieee_I1394 (.Y(N653), .A(inst_cellmath__7), .B(N652));
NOR3BXL inst_cellmath__70_0_I1395 (.Y(N5790), .AN(N653), .B(inst_cellmath__8), .C(inst_cellmath__4));
AND2X1 inst_cellmath__70_0_I1396 (.Y(inst_cellmath__70), .A(inst_cellmath__62), .B(N5790));
INVX2 inst_cellmath__73_0_I2603 (.Y(N7138), .A(N5751));
INVX3 inst_cellmath__73_0_I2608 (.Y(N7143), .A(N7138));
INVXL inst_cellmath__73_0_I2606 (.Y(N7141), .A(N7138));
INVXL inst_cellmath__73_0_I2605 (.Y(N7140), .A(N7138));
INVXL inst_cellmath__73_0_I2604 (.Y(N7139), .A(N7138));
NOR2X4 inst_cellmath__73_0_I1398 (.Y(N5875), .A(inst_cellmath__63), .B(N5751));
NOR2BX4 inst_cellmath__73_0_I1399 (.Y(N5820), .AN(inst_cellmath__63), .B(N7143));
AOI22XL inst_cellmath__73_0_I1400 (.Y(N5804), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[0]));
AOI22XL inst_cellmath__73_0_I1401 (.Y(N5847), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[1]));
AOI22XL inst_cellmath__73_0_I1402 (.Y(N5889), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[2]));
AOI22XL inst_cellmath__73_0_I1403 (.Y(N5834), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[3]));
AOI22XL inst_cellmath__73_0_I1404 (.Y(N5877), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[4]));
AOI22XL inst_cellmath__73_0_I1405 (.Y(N5821), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[5]));
AOI22XL inst_cellmath__73_0_I1406 (.Y(N5864), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[6]));
AOI22XL inst_cellmath__73_0_I1407 (.Y(N5808), .A0(inst_cellmath__70), .A1(N5875), .B0(N7143), .B1(inst_cellmath__57[7]));
AOI22XL inst_cellmath__73_0_I1408 (.Y(N5851), .A0(inst_cellmath__70), .A1(N5875), .B0(N7141), .B1(inst_cellmath__57[8]));
AOI22XL inst_cellmath__73_0_I1409 (.Y(N5796), .A0(inst_cellmath__70), .A1(N5875), .B0(N7141), .B1(inst_cellmath__57[9]));
AOI22XL inst_cellmath__73_0_I1410 (.Y(N5839), .A0(inst_cellmath__70), .A1(N5875), .B0(N7141), .B1(inst_cellmath__57[10]));
AOI22XL inst_cellmath__73_0_I1411 (.Y(N5881), .A0(inst_cellmath__70), .A1(N5875), .B0(N7141), .B1(inst_cellmath__57[11]));
AOI22XL inst_cellmath__73_0_I1412 (.Y(N5825), .A0(inst_cellmath__70), .A1(N5875), .B0(N7141), .B1(inst_cellmath__57[12]));
AOI22XL inst_cellmath__73_0_I1413 (.Y(N5868), .A0(inst_cellmath__70), .A1(N5875), .B0(N7140), .B1(inst_cellmath__57[13]));
AOI22XL inst_cellmath__73_0_I1414 (.Y(N5812), .A0(inst_cellmath__70), .A1(N5875), .B0(N7140), .B1(inst_cellmath__57[14]));
AOI22XL inst_cellmath__73_0_I1415 (.Y(N5856), .A0(inst_cellmath__70), .A1(N5875), .B0(N7140), .B1(inst_cellmath__57[15]));
AOI22XL inst_cellmath__73_0_I1416 (.Y(N5801), .A0(inst_cellmath__70), .A1(N5875), .B0(N7140), .B1(inst_cellmath__57[16]));
AOI22XL inst_cellmath__73_0_I1417 (.Y(N5844), .A0(inst_cellmath__70), .A1(N5875), .B0(N7140), .B1(inst_cellmath__57[17]));
AOI22XL inst_cellmath__73_0_I1418 (.Y(N5886), .A0(inst_cellmath__70), .A1(N5875), .B0(N7139), .B1(inst_cellmath__57[18]));
AOI22XL inst_cellmath__73_0_I1419 (.Y(N5831), .A0(inst_cellmath__70), .A1(N5875), .B0(N7139), .B1(inst_cellmath__57[19]));
AOI22XL inst_cellmath__73_0_I1420 (.Y(N5873), .A0(inst_cellmath__70), .A1(N5875), .B0(N7139), .B1(inst_cellmath__57[20]));
AOI22XL inst_cellmath__73_0_I1421 (.Y(N5817), .A0(inst_cellmath__70), .A1(N5875), .B0(N7139), .B1(inst_cellmath__57[21]));
AOI22XL inst_cellmath__73_0_I1422 (.Y(N5860), .A0(inst_cellmath__70), .A1(N5875), .B0(N7139), .B1(inst_cellmath__57[22]));
OAI2BB1XL inst_cellmath__73_0_I1423 (.Y(x[0]), .A0N(N5820), .A1N(inst_cellmath__64[0]), .B0(N5804));
OAI2BB1XL inst_cellmath__73_0_I1424 (.Y(x[1]), .A0N(N5820), .A1N(inst_cellmath__64[1]), .B0(N5847));
OAI2BB1XL inst_cellmath__73_0_I1425 (.Y(x[2]), .A0N(N5820), .A1N(inst_cellmath__64[2]), .B0(N5889));
OAI2BB1XL inst_cellmath__73_0_I1426 (.Y(x[3]), .A0N(N5820), .A1N(inst_cellmath__64[3]), .B0(N5834));
OAI2BB1XL inst_cellmath__73_0_I1427 (.Y(x[4]), .A0N(N5820), .A1N(inst_cellmath__64[4]), .B0(N5877));
OAI2BB1XL inst_cellmath__73_0_I1428 (.Y(x[5]), .A0N(N5820), .A1N(inst_cellmath__64[5]), .B0(N5821));
OAI2BB1XL inst_cellmath__73_0_I1429 (.Y(x[6]), .A0N(N5820), .A1N(inst_cellmath__64[6]), .B0(N5864));
OAI2BB1XL inst_cellmath__73_0_I1430 (.Y(x[7]), .A0N(N5820), .A1N(inst_cellmath__64[7]), .B0(N5808));
OAI2BB1XL inst_cellmath__73_0_I1431 (.Y(x[8]), .A0N(N5820), .A1N(inst_cellmath__64[8]), .B0(N5851));
OAI2BB1XL inst_cellmath__73_0_I1432 (.Y(x[9]), .A0N(N5820), .A1N(inst_cellmath__64[9]), .B0(N5796));
OAI2BB1XL inst_cellmath__73_0_I1433 (.Y(x[10]), .A0N(N5820), .A1N(inst_cellmath__64[10]), .B0(N5839));
OAI2BB1XL inst_cellmath__73_0_I1434 (.Y(x[11]), .A0N(N5820), .A1N(inst_cellmath__64[11]), .B0(N5881));
OAI2BB1XL inst_cellmath__73_0_I1435 (.Y(x[12]), .A0N(N5820), .A1N(inst_cellmath__64[12]), .B0(N5825));
OAI2BB1XL inst_cellmath__73_0_I1436 (.Y(x[13]), .A0N(N5820), .A1N(inst_cellmath__64[13]), .B0(N5868));
OAI2BB1XL inst_cellmath__73_0_I1437 (.Y(x[14]), .A0N(N5820), .A1N(inst_cellmath__64[14]), .B0(N5812));
OAI2BB1XL inst_cellmath__73_0_I1438 (.Y(x[15]), .A0N(N5820), .A1N(inst_cellmath__64[15]), .B0(N5856));
OAI2BB1XL inst_cellmath__73_0_I1439 (.Y(x[16]), .A0N(N5820), .A1N(inst_cellmath__64[16]), .B0(N5801));
OAI2BB1XL inst_cellmath__73_0_I1440 (.Y(x[17]), .A0N(N5820), .A1N(inst_cellmath__64[17]), .B0(N5844));
OAI2BB1XL inst_cellmath__73_0_I1441 (.Y(x[18]), .A0N(N5820), .A1N(inst_cellmath__64[18]), .B0(N5886));
OAI2BB1XL inst_cellmath__73_0_I1442 (.Y(x[19]), .A0N(N5820), .A1N(inst_cellmath__64[19]), .B0(N5831));
OAI2BB1XL inst_cellmath__73_0_I1443 (.Y(x[20]), .A0N(N5820), .A1N(inst_cellmath__64[20]), .B0(N5873));
OAI2BB1XL inst_cellmath__73_0_I1444 (.Y(x[21]), .A0N(N5820), .A1N(inst_cellmath__64[21]), .B0(N5817));
NAND2BXL inst_cellmath__73_0_I1445 (.Y(x[22]), .AN(N5820), .B(N5860));
assign inst_cellmath__27[0] = 1'B0;
assign inst_cellmath__33[0] = 1'B0;
assign inst_cellmath__33[1] = 1'B0;
assign inst_cellmath__33[2] = 1'B0;
assign inst_cellmath__33[3] = 1'B0;
assign inst_cellmath__33[4] = 1'B0;
assign inst_cellmath__33[5] = 1'B0;
assign inst_cellmath__33[6] = 1'B0;
assign inst_cellmath__33[7] = 1'B0;
assign inst_cellmath__33[8] = 1'B0;
assign inst_cellmath__33[9] = 1'B0;
assign inst_cellmath__33[10] = 1'B0;
assign inst_cellmath__33[11] = 1'B0;
assign inst_cellmath__33[12] = 1'B0;
assign inst_cellmath__33[13] = 1'B0;
assign inst_cellmath__33[14] = 1'B0;
assign inst_cellmath__33[15] = 1'B0;
assign inst_cellmath__33[16] = 1'B0;
assign inst_cellmath__33[17] = 1'B0;
assign inst_cellmath__33[18] = 1'B0;
assign inst_cellmath__33[19] = 1'B0;
assign inst_cellmath__33[20] = 1'B0;
assign inst_cellmath__33[21] = 1'B0;
assign inst_cellmath__33[22] = 1'B0;
assign inst_cellmath__33[23] = 1'B0;
assign inst_cellmath__33[29] = 1'B0;
assign inst_cellmath__33[31] = 1'B0;
assign inst_cellmath__33[33] = 1'B0;
assign inst_cellmath__33[35] = 1'B0;
assign inst_cellmath__33[37] = 1'B0;
assign inst_cellmath__33[39] = 1'B0;
assign inst_cellmath__35[0] = 1'B0;
assign inst_cellmath__36[0] = 1'B0;
assign inst_cellmath__36[1] = 1'B0;
assign inst_cellmath__36[2] = 1'B0;
assign inst_cellmath__36[3] = 1'B0;
assign inst_cellmath__36[4] = 1'B0;
assign inst_cellmath__36[5] = 1'B0;
assign inst_cellmath__36[6] = 1'B0;
assign inst_cellmath__36[7] = 1'B0;
assign inst_cellmath__36[8] = 1'B0;
assign inst_cellmath__36[9] = 1'B0;
assign inst_cellmath__36[10] = 1'B0;
assign inst_cellmath__36[11] = 1'B0;
assign inst_cellmath__36[12] = 1'B0;
assign inst_cellmath__36[13] = 1'B0;
assign inst_cellmath__36[14] = 1'B0;
assign inst_cellmath__36[15] = 1'B0;
assign inst_cellmath__36[16] = 1'B0;
assign inst_cellmath__36[17] = 1'B0;
assign inst_cellmath__36[18] = 1'B0;
assign inst_cellmath__36[19] = 1'B0;
assign inst_cellmath__36[20] = 1'B0;
assign inst_cellmath__36[21] = 1'B0;
assign inst_cellmath__36[22] = 1'B0;
assign inst_cellmath__36[23] = 1'B0;
assign inst_cellmath__36[24] = 1'B0;
assign inst_cellmath__36[25] = 1'B0;
assign inst_cellmath__36[49] = 1'B1;
assign inst_cellmath__37[11] = 1'B0;
assign inst_cellmath__37[13] = 1'B0;
assign inst_cellmath__37[14] = 1'B0;
assign inst_cellmath__37[15] = 1'B0;
assign inst_cellmath__37[16] = 1'B0;
assign inst_cellmath__37[18] = 1'B0;
assign inst_cellmath__37[20] = 1'B0;
assign inst_cellmath__37[21] = 1'B0;
assign inst_cellmath__37[22] = 1'B0;
assign inst_cellmath__37[23] = 1'B0;
assign inst_cellmath__37[42] = 1'B0;
assign inst_cellmath__37[43] = 1'B0;
assign inst_cellmath__37[44] = 1'B0;
assign inst_cellmath__37[45] = 1'B0;
assign inst_cellmath__37[46] = 1'B0;
assign inst_cellmath__37[47] = 1'B0;
assign inst_cellmath__37[48] = 1'B0;
assign inst_cellmath__37[49] = 1'B0;
assign inst_cellmath__45[26] = 1'B0;
assign inst_cellmath__49[0] = 1'B0;
assign inst_cellmath__49[2] = 1'B0;
assign inst_cellmath__49[3] = 1'B0;
assign inst_cellmath__50[0] = 1'B0;
assign inst_cellmath__59[8] = 1'B0;
assign inst_cellmath__59[9] = 1'B0;
assign inst_cellmath__64[22] = 1'B1;
assign inst_cellmath__68[1] = 1'B0;
assign inst_cellmath__68[2] = 1'B0;
assign inst_cellmath__68[3] = 1'B0;
assign inst_cellmath__68[4] = 1'B0;
assign inst_cellmath__68[5] = 1'B0;
assign inst_cellmath__68[6] = 1'B0;
assign inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  urH3Tw7Zoxg= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



