/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:00 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_2_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__9,
	inst_cellmath__17;
wire [8:0] inst_cellmath__19;
wire [7:0] inst_cellmath__20;
wire [8:0] inst_cellmath__22;
wire  inst_cellmath__29,
	inst_cellmath__33,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42;
wire [18:0] inst_cellmath__51;
wire [39:0] inst_cellmath__62__W0, inst_cellmath__62__W1,
	inst_cellmath__63__W0, inst_cellmath__63__W1;
wire [39:0] inst_cellmath__64;
wire  inst_cellmath__67;
wire N446,N447,N448,N449,N450,N451,N452 
	,N453,N454,N455,N456,N457,N477,N478,N479 
	,N480,N481,N482,N483,N484,N485,N486,N487 
	,N488,N489,N490,N491,N492,N493,N494,N495 
	,N496,N497,N498,N499,N500,N2353,N2355,N2376 
	,N2378,N2381,N2384,N2387,N2389,N2393,N2395,N2402 
	,N2404,N2408,N2444,N2449,N2451,N2454,N2457,N2459 
	,N2464,N2483,N2486,N2489,N2514,N2516,N2518,N2523 
	,N2526,N2576,N2577,N2578,N2579,N2580,N2581,N2583 
	,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591 
	,N2592,N2593,N2595,N2596,N2597,N2599,N2600,N2601 
	,N2602,N2603,N2604,N2605,N2606,N2608,N2609,N2610 
	,N2611,N2614,N2615,N2616,N2617,N2619,N2620,N2621 
	,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630 
	,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638 
	,N2639,N2641,N2642,N2643,N2644,N2645,N2647,N2648 
	,N2649,N2650,N2652,N2655,N2656,N2658,N2659,N2660 
	,N2661,N2663,N2665,N2666,N2667,N2668,N2670,N2671 
	,N2672,N2673,N2674,N2675,N2677,N2678,N2679,N2680 
	,N2681,N2682,N2683,N2684,N2685,N2686,N2688,N2689 
	,N2690,N2691,N2694,N2695,N2696,N2697,N2698,N2699 
	,N2701,N2702,N2703,N2704,N2705,N2706,N2708,N2709 
	,N2710,N2711,N2712,N2713,N2714,N2715,N2717,N2719 
	,N2720,N2721,N2722,N2723,N2724,N2726,N2727,N2729 
	,N2730,N2731,N2732,N2733,N2734,N2735,N2737,N2738 
	,N2740,N2741,N2742,N2744,N2745,N2746,N2747,N2748 
	,N2749,N2751,N2752,N2753,N2754,N2757,N2759,N2761 
	,N2762,N2763,N2765,N2766,N2767,N2768,N2769,N2770 
	,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778 
	,N2779,N2781,N2782,N2783,N2784,N2786,N2787,N2788 
	,N2789,N2790,N2791,N2793,N2794,N2796,N2797,N2798 
	,N2799,N2800,N2801,N2802,N2803,N2805,N2806,N2807 
	,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815 
	,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823 
	,N2824,N2826,N2827,N2828,N2829,N2830,N2831,N2832 
	,N2833,N2834,N2836,N2837,N2838,N2839,N2840,N2841 
	,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2850 
	,N2851,N2852,N2853,N2854,N2855,N2857,N2858,N2860 
	,N2861,N2862,N2864,N2865,N2867,N2868,N2869,N2870 
	,N2871,N2874,N2875,N2877,N2878,N2879,N2880,N2881 
	,N2883,N2884,N2885,N2886,N2887,N2888,N2890,N2891 
	,N2892,N2893,N2894,N2895,N3203,N3204,N3205,N3206 
	,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214 
	,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223 
	,N3224,N3225,N3226,N3227,N3229,N3230,N3231,N3232 
	,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240 
	,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248 
	,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257 
	,N3258,N3259,N3260,N3262,N3263,N3264,N3265,N3266 
	,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274 
	,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282 
	,N3283,N3285,N3286,N3287,N3288,N3289,N3290,N3291 
	,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299 
	,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308 
	,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316 
	,N3317,N3318,N3320,N3321,N3322,N3323,N3324,N3325 
	,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333 
	,N3334,N3335,N3336,N3338,N3339,N3340,N3341,N3342 
	,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350 
	,N3352,N3353,N3354,N3355,N3356,N3357,N3358,N3359 
	,N3360,N3361,N3362,N3363,N3364,N3365,N3367,N3368 
	,N3369,N3370,N3371,N3372,N3374,N3375,N3376,N3377 
	,N3378,N3379,N3380,N3381,N3382,N3383,N3385,N3386 
	,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394 
	,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402 
	,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410 
	,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3419 
	,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427 
	,N3428,N3429,N3430,N3431,N3432,N3434,N3435,N3436 
	,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444 
	,N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452 
	,N3453,N3455,N3456,N3457,N3458,N3459,N3460,N3461 
	,N3462,N3463,N3464,N3465,N3466,N3467,N3469,N3470 
	,N3471,N3472,N3473,N3474,N3475,N3476,N3477,N3478 
	,N3479,N3480,N3481,N3483,N3484,N3485,N3486,N3487 
	,N3488,N3489,N3490,N3491,N3492,N3494,N3495,N3496 
	,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504 
	,N3505,N3506,N3508,N3509,N3510,N3511,N3512,N3513 
	,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521 
	,N3522,N3523,N3524,N3526,N3527,N3528,N3529,N3530 
	,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538 
	,N3539,N3540,N3541,N3543,N3544,N3545,N3546,N3547 
	,N3548,N3549,N3550,N3551,N3553,N3554,N3555,N3556 
	,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564 
	,N3565,N3566,N3567,N3568,N3569,N3570,N3571,N3572 
	,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581 
	,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3590 
	,N3591,N3592,N3593,N3594,N3595,N3596,N3597,N3598 
	,N3599,N3600,N3601,N3603,N3604,N3605,N3606,N3607 
	,N3608,N3609,N3610,N3611,N3612,N3614,N3615,N3616 
	,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624 
	,N3625,N3626,N3627,N3629,N3630,N3631,N3632,N3633 
	,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641 
	,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650 
	,N3651,N3652,N3653,N3654,N3655,N3656,N3658,N3659 
	,N3660,N3661,N3662,N3663,N3664,N3666,N3667,N3668 
	,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3677 
	,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685 
	,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693 
	,N3694,N3695,N3697,N3698,N3699,N3700,N3701,N3702 
	,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3711 
	,N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719 
	,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727 
	,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736 
	,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744 
	,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753 
	,N3754,N3755,N3756,N3757,N3758,N3759,N3761,N3762 
	,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770 
	,N3771,N3773,N3774,N3775,N3776,N3777,N3779,N3780 
	,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788 
	,N3789,N3790,N3791,N3792,N3793,N3794,N3796,N3797 
	,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805 
	,N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813 
	,N3814,N3816,N3817,N3818,N3819,N3820,N3821,N3822 
	,N3823,N3824,N3825,N3826,N3827,N3828,N3830,N3831 
	,N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839 
	,N3840,N3842,N3843,N3844,N3845,N3846,N3847,N3848 
	,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857 
	,N3858,N3859,N3860,N3861,N3862,N3864,N3865,N3866 
	,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874 
	,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883 
	,N3884,N3885,N3886,N3887,N3889,N3890,N3891,N3892 
	,N3893,N3894,N3895,N3896,N3897,N3899,N3900,N3901 
	,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909 
	,N3910,N3911,N3912,N3913,N3915,N3916,N3917,N3918 
	,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926 
	,N3927,N3928,N3929,N3930,N3931,N3933,N3934,N3935 
	,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943 
	,N3944,N3945,N3946,N3947,N3949,N3950,N3951,N3952 
	,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3962 
	,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970 
	,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3979 
	,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987 
	,N3988,N3989,N3990,N3992,N3993,N3994,N3995,N3996 
	,N3997,N3998,N3999,N4000,N4001,N4002,N4004,N4005 
	,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013 
	,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022 
	,N4023,N4024,N4025,N4027,N4028,N4029,N4030,N4031 
	,N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039 
	,N4040,N4041,N4042,N4043,N4044,N4046,N4047,N4048 
	,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056 
	,N4057,N4059,N4060,N4061,N4062,N4063,N4065,N4066 
	,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074 
	,N4075,N4076,N4077,N4078,N4079,N4080,N4082,N4083 
	,N4084,N4085,N4086,N4087,N4088,N4089,N4090,N4091 
	,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099 
	,N4100,N4101,N4102,N4103,N4104,N4106,N4107,N4108 
	,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116 
	,N4117,N4118,N4120,N4121,N4122,N4123,N4124,N4125 
	,N4126,N4127,N4128,N4130,N4131,N4132,N4133,N4134 
	,N4135,N5062,N5064,N5066,N5067,N5069,N5070,N5071 
	,N5072,N5073,N5075,N5076,N5077,N5078,N5079,N5080 
	,N5081,N5083,N5084,N5085,N5086,N5087,N5088,N5089 
	,N5090,N5091,N5092,N5094,N5095,N5097,N5098,N5099 
	,N5101,N5102,N5104,N5105,N5106,N5108,N5110,N5111 
	,N5112,N5113,N5114,N5115,N5116,N5118,N5119,N5120 
	,N5121,N5122,N5123,N5125,N5126,N5127,N5129,N5130 
	,N5131,N5132,N5133,N5134,N5135,N5137,N5138,N5139 
	,N5141,N5143,N5144,N5145,N5146,N5147,N5148,N5150 
	,N5151,N5152,N5153,N5154,N5155,N5156,N5157,N5158 
	,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5169 
	,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178 
	,N5179,N5182,N5183,N5184,N5185,N5186,N5187,N5189 
	,N5190,N5192,N5193,N5194,N5195,N5196,N5197,N5198 
	,N5199,N5201,N5203,N5204,N5205,N5206,N5207,N5208 
	,N5209,N5211,N5212,N5214,N5215,N5216,N5217,N5218 
	,N5219,N5220,N5221,N5223,N5224,N5226,N5228,N5229 
	,N5231,N5232,N5233,N5234,N5235,N5236,N5237,N5238 
	,N5240,N5241,N5242,N5244,N5245,N5246,N5247,N5248 
	,N5249,N5250,N5252,N5254,N5255,N5256,N5257,N5258 
	,N5259,N5260,N5261,N5263,N5264,N5265,N5266,N5267 
	,N5268,N5269,N5270,N5272,N5273,N5274,N5276,N5277 
	,N5278,N5279,N5280,N5281,N5283,N5284,N5286,N5287 
	,N5289,N5290,N5291,N5292,N5293,N5295,N5296,N5297 
	,N5299,N5300,N5301,N5302,N5303,N5304,N5305,N5307 
	,N5308,N5309,N5310,N5311,N5312,N5313,N5315,N5316 
	,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325 
	,N5326,N5327,N5328,N5330,N5332,N5333,N5334,N5335 
	,N5337,N5338,N5339,N5340,N5341,N5342,N5343,N5344 
	,N5345,N5346,N5347,N5349,N5352,N5353,N5354,N5355 
	,N5356,N5357,N5358,N5361,N5362,N5363,N5364,N5365 
	,N5366,N5367,N5368,N5370,N5371,N5372,N5374,N5376 
	,N5377,N5378,N5379,N5380,N5381,N5382,N5384,N5385 
	,N5386,N5387,N5388,N5389,N5390,N5391,N5393,N5395 
	,N5396,N5397,N5398,N5399,N5400,N5401,N5721,N5722 
	,N5723,N5724,N5726,N5728,N5729,N5730,N5731,N5732 
	,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740 
	,N5741,N5742,N5743,N5744,N5745,N5747,N5748,N5749 
	,N5751,N5752,N5753,N5754,N5756,N5757,N5758,N5759 
	,N5760,N5762,N5763,N5764,N5765,N5766,N5767,N5769 
	,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777 
	,N5778,N5779,N5780,N5782,N5783,N5784,N5785,N5787 
	,N5788,N5789,N5790,N5791,N5792,N5793,N5795,N5796 
	,N5797,N5798,N5799,N5800,N5801,N5802,N5804,N5805 
	,N5806,N5807,N5808,N5809,N5810,N5811,N5812,N5813 
	,N5814,N5816,N5818,N5819,N5820,N5821,N5822,N5823 
	,N5824,N5825,N5827,N5828,N5829,N5831,N5832,N5833 
	,N5834,N5836,N5837,N5838,N5839,N5840,N5841,N5842 
	,N5844,N5845,N5846,N5847,N5848,N5849,N5850,N5851 
	,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859 
	,N5861,N5862,N5863,N5864,N5865,N5867,N5868,N5870 
	,N5871,N5872,N5873,N5874,N5875,N5877,N5878,N5879 
	,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887 
	,N5888,N5889,N5890,N5892,N5893,N5894,N5895,N5896 
	,N5897,N5898,N5899,N5901,N5902,N5903,N5904,N5905 
	,N5906,N5909,N5910,N5912,N5913,N5914,N5915,N5916 
	,N5917,N5918,N5919,N5920,N5921,N5922,N5925,N5926 
	,N5927,N5928,N5929,N5930,N5931,N5932,N5933,N5935 
	,N5936,N5937,N5938,N5939,N5941,N5942,N5944,N5945 
	,N5946,N5947,N5948,N5949,N5950,N5952,N5953,N5954 
	,N5955,N5956,N5958,N5959,N5960,N5961,N5962,N5963 
	,N5964,N5965,N5966,N5967,N5968,N5969,N5970,N5971 
	,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980 
	,N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988 
	,N5990,N5991,N5992,N5993,N5994,N5995,N5996,N5997 
	,N5998,N5999,N6000,N6001,N6002,N6003,N6005,N6007 
	,N6008,N6009,N6010,N6011,N6012,N6014,N6015,N6016 
	,N6017,N6019,N6020,N6021,N6022,N6024,N6025,N6026 
	,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034 
	,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6044 
	,N6045,N6046,N6047,N6049,N6050,N6051,N6053,N6054 
	,N6055,N6056,N6058,N6059,N6060,N6061,N6062,N6063 
	,N6064,N6065,N6067,N6068,N6069,N6070,N6071,N6072 
	,N6073,N6074,N6075,N6076,N6077,N6078,N6079,N6080 
	,N6082,N6083,N6084,N6085,N6086,N6087,N6089,N6090 
	,N6091,N6093,N6094,N6095,N6096,N6098,N6099,N6100 
	,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6109 
	,N6110,N6113,N6114,N6115,N6116,N6117,N6118,N6119 
	,N6120,N6121,N6122,N6124,N6125,N6126,N6128,N6129 
	,N6130,N6131,N6132,N6134,N6135,N6136,N6137,N6138 
	,N6139,N6140,N6141,N6143,N6144,N6145,N6146,N6147 
	,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155 
	,N6156,N6158,N6159,N6160,N6161,N6162,N6163,N6165 
	,N6166,N6167,N6168,N6169,N6170,N6171,N6172,N6174 
	,N6175,N6177,N6178,N6179,N6180,N6181,N6182,N6183 
	,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6192 
	,N6193,N6194,N6195,N6196,N6197,N6198,N6199,N6201 
	,N6202,N6203,N6204,N6206,N6207,N6209,N6210,N6211 
	,N6212,N6213,N6214,N6215,N6216,N6217,N6218,N6220 
	,N6221,N6222,N6223,N6224,N6225,N6226,N6227,N6228 
	,N6230,N6231,N6232,N6233,N6234,N6237,N6238,N6240 
	,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248 
	,N6249,N6250,N6251,N6253,N6254,N6255,N6256,N6257 
	,N6258,N6259,N6260,N6261,N6262,N6263,N6264,N6265 
	,N6266,N6267,N6268,N6270,N6271,N6273,N6274,N6275 
	,N6276,N6278,N6279,N6280,N6281,N6282,N6283,N6284 
	,N6285,N6287,N6288,N6289,N6290,N6291,N6292,N6293 
	,N6294,N6295,N6296,N6297,N6299,N6300,N6301,N6302 
	,N6303,N6304,N6305,N6306,N6307,N6308,N6309,N6310 
	,N6313,N6314,N6315,N6316,N6318,N6319,N6320,N6322 
	,N6323,N6324,N6325,N6326,N6327,N6329,N6330,N6331 
	,N6332,N6333,N6335,N6336,N6337,N6338,N6339,N6340 
	,N6341,N6342,N6343,N6344,N6345,N6346,N6347,N6348 
	,N6350,N6351,N6352,N6354,N6355,N6356,N6357,N6358 
	,N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6367 
	,N6368,N6369,N6370,N6371,N6372,N6373,N6374,N6375 
	,N6376,N6377,N6378,N6380,N6381,N6382,N6384,N6385 
	,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6394 
	,N6395,N6396,N6398,N6399,N6401,N6402,N6403,N6404 
	,N6405,N6406,N6407,N6408,N6410,N6411,N6412,N6413 
	,N6414,N6415,N6416,N6417,N6418,N6419,N6420,N6422 
	,N6423,N6425,N6426,N6427,N6428,N6430,N6431,N6432 
	,N6433,N6434,N6435,N6436,N6437,N6439,N6440,N6442 
	,N6443,N6444,N6445,N6446,N6447,N6448,N6449,N6450 
	,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6459 
	,N6460,N6461,N6462,N6463,N6465,N6466,N6467,N6469 
	,N6470,N6471,N6472,N6473,N6474,N6475,N6477,N6478 
	,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486 
	,N6487,N6488,N6490,N6491,N6492,N6493,N6494,N6495 
	,N6496,N6498,N6499,N6500,N6501,N6502,N6503,N6506 
	,N6507,N6509,N6510,N6511,N6512,N6513,N6514,N6515 
	,N6516,N6517,N6519,N6520,N6521,N6522,N6523,N6524 
	,N6525,N6526,N6527,N6528,N6529,N6530,N6531,N6532 
	,N6533,N6534,N6535,N6536,N6537,N6538,N6540,N6541 
	,N6543,N6544,N6545,N6546,N6547,N6548,N6549,N6550 
	,N6551,N6552,N6553,N6555,N6556,N6557,N6558,N6559 
	,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6568 
	,N6569,N6570,N6572,N6573,N6574,N6575,N6576,N6577 
	,N6578,N6579,N7408,N7412,N7414,N7415,N7416,N7420 
	,N7423,N7427,N7431,N7432,N7436,N7438,N7440,N7442 
	,N7444,N7445,N7450,N7452,N7453,N7456,N7459,N7461 
	,N7465,N7467,N7468,N7474,N7476,N7477,N7478,N7479 
	,N7481,N7484,N7486,N7487,N7489,N7491,N7492,N7495 
	,N7500,N7503,N7505,N7506,N7510,N7512,N7514,N7515 
	,N7517,N7523,N7525,N7526,N7528,N7532,N7534,N7540 
	,N7543,N7544,N7546,N7547,N7548,N7549,N7550,N7551 
	,N7552,N7554,N7555,N7556,N7558,N7561,N7564,N7566 
	,N7568,N7570,N7571,N7572,N7574,N7579,N7581,N7583 
	,N7585,N7586,N7590,N7592,N7593,N7595,N7597,N7599 
	,N7602,N7604,N7605,N7607,N7609,N7612,N7614,N7617 
	,N7618,N7619,N7620,N7623,N7624,N7625,N7628,N7631 
	,N7634,N7636,N7637,N7639,N7641,N7642,N7647,N7651 
	,N7652,N7654,N7656,N7662,N7663,N7665,N7667,N7668 
	,N7669,N7673,N7676,N7678,N7686,N7688,N7689,N7690 
	,N7692,N7693,N7694,N7696,N7698,N7701,N7703,N7709 
	,N7711,N7713,N7715,N7716,N7720,N7722,N7723,N7730 
	,N7733,N7734,N7736,N7737,N7739,N7741,N7742,N7745 
	,N7753,N7755,N7757,N7758,N7762,N7763,N7764,N7765 
	,N7767,N7768,N7769,N7770,N7773,N7775,N7776,N7778 
	,N7779,N7783,N7785,N7786,N7787,N7789,N7790,N7791 
	,N7795,N7796,N7798,N7800,N7804,N7806,N7808,N7809 
	,N7811,N7812,N7814,N7817,N7819,N7823,N7825,N7827 
	,N7828,N7831,N7835,N7839,N7843,N7846,N7848,N7850 
	,N7851,N7852,N7853,N7854,N7857,N7859,N7860,N7861 
	,N7865,N7868,N7871,N7873,N7876,N7878,N7881,N7882 
	,N7886,N7887,N7889,N7891,N7893,N7895,N7902,N7903 
	,N7905,N7909,N7911,N7912,N7921,N7922,N7924,N7925 
	,N7926,N7927,N7929,N7931,N7933,N7934,N7940,N7943 
	,N7945,N7946,N7948,N7949,N7951,N7954,N7959,N7961 
	,N7962,N7963,N7964,N7967,N7969,N7970,N7971,N7972 
	,N7974,N7978,N7979,N7980,N7982,N7984,N7987,N7988 
	,N7990,N7991,N7992,N7993,N7995,N7996,N7997,N8001 
	,N8002,N8004,N8005,N11575,N11605,N22792,N22794,N22796 
	;
NAND2XL inst_cellmath__9_0_I160 (.Y(N2353), .A(a_exp[7]), .B(a_exp[0]));
AND4XL inst_cellmath__9_0_I13847 (.Y(N2355), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL hyperpropagate_4_1_A_I4939 (.Y(N11575), .A(a_exp[6]), .B(a_exp[5]), .C(N2355));
NOR2XL hyperpropagate_4_1_A_I4940 (.Y(inst_cellmath__9), .A(N2353), .B(N11575));
NOR2XL inst_cellmath__15__5__I169 (.Y(N2381), .A(a_man[18]), .B(a_man[17]));
NOR2XL inst_cellmath__15__5__I173 (.Y(N2376), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__15__5__I174 (.Y(N2384), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__15__5__I175 (.Y(N2395), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__15__5__I176 (.Y(N2404), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__15__5__I13848 (.Y(N2389), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__15__5__I13849 (.Y(N2408), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 inst_cellmath__15__5__I13850 (.Y(N2402), .AN(N2381), .B(a_man[16]), .C(N2408), .D(a_man[15]));
NOR4X1 inst_cellmath__15__5__I180 (.Y(N2393), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N2389));
NAND4XL inst_cellmath__15__5__I182 (.Y(N2387), .A(N2376), .B(N2395), .C(N2384), .D(N2404));
NAND2XL inst_cellmath__15__5__I183 (.Y(N2378), .A(N2393), .B(N2402));
NOR2XL inst_cellmath__15__5__I184 (.Y(inst_cellmath__19[0]), .A(N2387), .B(N2378));
NOR2BX1 cynw_cm_float_rcp_I185 (.Y(inst_cellmath__29), .AN(inst_cellmath__9), .B(inst_cellmath__19[0]));
NOR2BX1 cynw_cm_float_rcp_I186 (.Y(x[31]), .AN(a_sign), .B(inst_cellmath__29));
INVXL cynw_cm_float_rcp_I5 (.Y(inst_cellmath__20[0]), .A(a_exp[0]));
INVXL cynw_cm_float_rcp_I6 (.Y(inst_cellmath__20[1]), .A(a_exp[1]));
INVXL cynw_cm_float_rcp_I8 (.Y(inst_cellmath__20[3]), .A(a_exp[3]));
INVXL cynw_cm_float_rcp_I10 (.Y(inst_cellmath__20[5]), .A(a_exp[5]));
INVXL cynw_cm_float_rcp_I12 (.Y(inst_cellmath__20[7]), .A(a_exp[7]));
ADDHX1 inst_cellmath__22_0_I188 (.CO(N2464), .S(inst_cellmath__22[0]), .A(inst_cellmath__20[0]), .B(inst_cellmath__19[0]));
XNOR2X1 inst_cellmath__22_0_I189 (.Y(inst_cellmath__22[1]), .A(inst_cellmath__20[1]), .B(N2464));
NOR2XL inst_cellmath__22_0_I190 (.Y(N2459), .A(inst_cellmath__20[1]), .B(N2464));
XNOR2X1 inst_cellmath__22_0_I191 (.Y(inst_cellmath__22[2]), .A(a_exp[2]), .B(N2459));
NAND2XL inst_cellmath__22_0_I192 (.Y(N2457), .A(a_exp[2]), .B(N2459));
XNOR2X1 inst_cellmath__22_0_I193 (.Y(inst_cellmath__22[3]), .A(inst_cellmath__20[3]), .B(N2457));
NOR2XL inst_cellmath__22_0_I194 (.Y(N2454), .A(inst_cellmath__20[3]), .B(N2457));
XNOR2X1 inst_cellmath__22_0_I195 (.Y(inst_cellmath__22[4]), .A(a_exp[4]), .B(N2454));
NAND2XL inst_cellmath__22_0_I196 (.Y(N2451), .A(a_exp[4]), .B(N2454));
XNOR2X1 inst_cellmath__22_0_I197 (.Y(inst_cellmath__22[5]), .A(inst_cellmath__20[5]), .B(N2451));
NOR2XL inst_cellmath__22_0_I198 (.Y(N2449), .A(inst_cellmath__20[5]), .B(N2451));
XNOR2X1 inst_cellmath__22_0_I199 (.Y(inst_cellmath__22[6]), .A(a_exp[6]), .B(N2449));
NAND2XL inst_cellmath__22_0_I200 (.Y(N2444), .A(a_exp[6]), .B(N2449));
XNOR2X1 inst_cellmath__22_0_I201 (.Y(inst_cellmath__22[7]), .A(inst_cellmath__20[7]), .B(N2444));
NOR3XL inst_cellmath__17__6__I203 (.Y(N2486), .A(inst_cellmath__22[2]), .B(inst_cellmath__22[3]), .C(inst_cellmath__22[5]));
NOR2XL inst_cellmath__17__6__I204 (.Y(N2489), .A(inst_cellmath__22[6]), .B(inst_cellmath__22[7]));
NOR4BX1 inst_cellmath__17__6__I205 (.Y(N2483), .AN(N2489), .B(inst_cellmath__22[0]), .C(inst_cellmath__22[4]), .D(inst_cellmath__22[1]));
NAND2XL inst_cellmath__17__6__I206 (.Y(N446), .A(N2486), .B(N2483));
OAI21XL cynw_cm_float_rcp_I4901 (.Y(inst_cellmath__17), .A0(inst_cellmath__20[7]), .A1(N2444), .B0(N446));
MX2XL cynw_cm_float_rcp_I4933 (.Y(N447), .A(inst_cellmath__17), .B(inst_cellmath__19[0]), .S0(inst_cellmath__9));
NOR2BX1 cynw_cm_float_rcp_I210 (.Y(inst_cellmath__33), .AN(N447), .B(inst_cellmath__29));
NOR2XL inst_cellmath__34_0_I211 (.Y(N2523), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL inst_cellmath__34_0_I212 (.Y(N2526), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL inst_cellmath__34_0_I213 (.Y(N2514), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL inst_cellmath__34_0_I214 (.Y(N2518), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL inst_cellmath__34_0_I215 (.Y(N2516), .A(N2523), .B(N2514), .C(N2526), .D(N2518));
NOR2XL inst_cellmath__34_0_I216 (.Y(inst_cellmath__34), .A(N2516), .B(inst_cellmath__29));
NOR3XL cynw_cm_float_rcp_I217 (.Y(inst_cellmath__42), .A(inst_cellmath__29), .B(inst_cellmath__34), .C(inst_cellmath__33));
OR2XL cynw_cm_float_rcp_I218 (.Y(inst_cellmath__38), .A(inst_cellmath__29), .B(inst_cellmath__34));
MX2XL inst_cellmath__43_0_I219 (.Y(x[23]), .A(inst_cellmath__38), .B(inst_cellmath__22[0]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I220 (.Y(x[24]), .A(inst_cellmath__38), .B(inst_cellmath__22[1]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I221 (.Y(x[25]), .A(inst_cellmath__38), .B(inst_cellmath__22[2]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I222 (.Y(x[26]), .A(inst_cellmath__38), .B(inst_cellmath__22[3]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I223 (.Y(x[27]), .A(inst_cellmath__38), .B(inst_cellmath__22[4]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I224 (.Y(x[28]), .A(inst_cellmath__38), .B(inst_cellmath__22[5]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I225 (.Y(x[29]), .A(inst_cellmath__38), .B(inst_cellmath__22[6]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I226 (.Y(x[30]), .A(inst_cellmath__38), .B(inst_cellmath__22[7]), .S0(inst_cellmath__42));
OR4X1 cynw_cm_float_rcp_I227 (.Y(N448), .A(inst_cellmath__19[0]), .B(inst_cellmath__29), .C(inst_cellmath__34), .D(inst_cellmath__33));
INVXL cynw_cm_float_rcp_I24 (.Y(inst_cellmath__67), .A(N448));
INVXL cynw_cm_float_rcp_I25 (.Y(inst_cellmath__63__W0[33]), .A(a_man[15]));
INVXL inst_cellmath__60_0_I228 (.Y(N2631), .A(a_man[4]));
INVXL inst_cellmath__60_0_I229 (.Y(N2698), .A(a_man[5]));
INVXL inst_cellmath__60_0_I230 (.Y(N2772), .A(a_man[6]));
INVXL inst_cellmath__60_0_I231 (.Y(N2579), .A(a_man[7]));
INVXL inst_cellmath__60_0_I232 (.Y(N2648), .A(a_man[8]));
INVXL inst_cellmath__60_0_I233 (.Y(N2746), .A(a_man[9]));
INVXL inst_cellmath__60_0_I234 (.Y(N2822), .A(a_man[10]));
INVXL inst_cellmath__60_0_I235 (.Y(N2887), .A(a_man[11]));
INVXL inst_cellmath__60_0_I236 (.Y(N2637), .A(a_man[12]));
INVXL inst_cellmath__60_0_I237 (.Y(N2705), .A(a_man[13]));
INVXL inst_cellmath__60_0_I238 (.Y(N2776), .A(a_man[14]));
INVXL inst_cellmath__60_0_I239 (.Y(N2847), .A(inst_cellmath__63__W0[33]));
INVXL inst_cellmath__60_0_I240 (.Y(N2875), .A(a_man[3]));
NOR2XL inst_cellmath__60_0_I243 (.Y(N2675), .A(N2875), .B(N2772));
NOR2XL inst_cellmath__60_0_I244 (.Y(N2821), .A(N2875), .B(N2579));
NOR2XL inst_cellmath__60_0_I245 (.Y(N2636), .A(N2875), .B(N2648));
NOR2XL inst_cellmath__60_0_I246 (.Y(N2778), .A(N2875), .B(N2746));
NOR2XL inst_cellmath__60_0_I247 (.Y(N2595), .A(N2875), .B(N2822));
NOR2XL inst_cellmath__60_0_I248 (.Y(N2732), .A(N2875), .B(N2887));
NOR2XL inst_cellmath__60_0_I249 (.Y(N2877), .A(N2875), .B(N2637));
NOR2XL inst_cellmath__60_0_I250 (.Y(N2691), .A(N2875), .B(N2705));
NOR2XL inst_cellmath__60_0_I251 (.Y(N2838), .A(N2875), .B(N2776));
OR2XL inst_cellmath__60_0_I252 (.Y(N2611), .A(N2875), .B(N2847));
NOR2XL inst_cellmath__60_0_I253 (.Y(N2814), .A(N2631), .B(N2698));
NOR2XL inst_cellmath__60_0_I254 (.Y(N2629), .A(N2631), .B(N2772));
NOR2XL inst_cellmath__60_0_I255 (.Y(N2770), .A(N2631), .B(N2579));
NOR2XL inst_cellmath__60_0_I256 (.Y(N2590), .A(N2631), .B(N2648));
NOR2XL inst_cellmath__60_0_I257 (.Y(N2727), .A(N2631), .B(N2746));
NOR2XL inst_cellmath__60_0_I258 (.Y(N2867), .A(N2631), .B(N2822));
NOR2XL inst_cellmath__60_0_I259 (.Y(N2685), .A(N2631), .B(N2887));
NOR2XL inst_cellmath__60_0_I260 (.Y(N2833), .A(N2631), .B(N2637));
NOR2XL inst_cellmath__60_0_I261 (.Y(N2647), .A(N2631), .B(N2705));
NOR2XL inst_cellmath__60_0_I262 (.Y(N2789), .A(N2631), .B(N2776));
OR2XL inst_cellmath__60_0_I263 (.Y(N2679), .A(N2631), .B(N2847));
INVXL inst_cellmath__60_0_I264 (.Y(N2807), .A(N2698));
NOR2XL inst_cellmath__60_0_I265 (.Y(N2762), .A(N2698), .B(N2772));
NOR2XL inst_cellmath__60_0_I266 (.Y(N2585), .A(N2698), .B(N2579));
NOR2XL inst_cellmath__60_0_I267 (.Y(N2721), .A(N2698), .B(N2648));
NOR2XL inst_cellmath__60_0_I268 (.Y(N2861), .A(N2698), .B(N2746));
NOR2XL inst_cellmath__60_0_I269 (.Y(N2680), .A(N2698), .B(N2822));
NOR2XL inst_cellmath__60_0_I270 (.Y(N2829), .A(N2698), .B(N2887));
NOR2XL inst_cellmath__60_0_I271 (.Y(N2643), .A(N2698), .B(N2637));
NOR2XL inst_cellmath__60_0_I272 (.Y(N2784), .A(N2698), .B(N2705));
NOR2XL inst_cellmath__60_0_I273 (.Y(N2602), .A(N2698), .B(N2776));
OR2XL inst_cellmath__60_0_I274 (.Y(N2752), .A(N2698), .B(N2847));
INVXL inst_cellmath__60_0_I275 (.Y(N2616), .A(N2772));
NOR2XL inst_cellmath__60_0_I276 (.Y(N2578), .A(N2772), .B(N2579));
NOR2XL inst_cellmath__60_0_I277 (.Y(N2715), .A(N2772), .B(N2648));
NOR2XL inst_cellmath__60_0_I278 (.Y(N2855), .A(N2772), .B(N2746));
NOR2XL inst_cellmath__60_0_I279 (.Y(N2673), .A(N2772), .B(N2822));
NOR2XL inst_cellmath__60_0_I280 (.Y(N2819), .A(N2772), .B(N2887));
NOR2XL inst_cellmath__60_0_I281 (.Y(N2635), .A(N2772), .B(N2637));
NOR2XL inst_cellmath__60_0_I282 (.Y(N2775), .A(N2772), .B(N2705));
NOR2XL inst_cellmath__60_0_I283 (.Y(N2593), .A(N2772), .B(N2776));
OR2XL inst_cellmath__60_0_I284 (.Y(N2828), .A(N2772), .B(N2847));
INVXL inst_cellmath__60_0_I285 (.Y(N2609), .A(N2579));
NOR2XL inst_cellmath__60_0_I286 (.Y(N2891), .A(N2579), .B(N2648));
NOR2XL inst_cellmath__60_0_I287 (.Y(N2709), .A(N2579), .B(N2746));
NOR2XL inst_cellmath__60_0_I288 (.Y(N2850), .A(N2579), .B(N2822));
NOR2XL inst_cellmath__60_0_I289 (.Y(N2666), .A(N2579), .B(N2887));
NOR2XL inst_cellmath__60_0_I290 (.Y(N2811), .A(N2579), .B(N2637));
NOR2XL inst_cellmath__60_0_I291 (.Y(N2624), .A(N2579), .B(N2705));
NOR2XL inst_cellmath__60_0_I292 (.Y(N2767), .A(N2579), .B(N2776));
OR2XL inst_cellmath__60_0_I293 (.Y(N2893), .A(N2579), .B(N2847));
INVXL inst_cellmath__60_0_I294 (.Y(N2787), .A(N2648));
NOR2XL inst_cellmath__60_0_I295 (.Y(N2741), .A(N2648), .B(N2746));
NOR2XL inst_cellmath__60_0_I296 (.Y(N2884), .A(N2648), .B(N2822));
NOR2XL inst_cellmath__60_0_I297 (.Y(N2701), .A(N2648), .B(N2887));
NOR2XL inst_cellmath__60_0_I298 (.Y(N2844), .A(N2648), .B(N2637));
NOR2XL inst_cellmath__60_0_I299 (.Y(N2659), .A(N2648), .B(N2705));
NOR2XL inst_cellmath__60_0_I300 (.Y(N2803), .A(N2648), .B(N2776));
OR2XL inst_cellmath__60_0_I301 (.Y(N2642), .A(N2648), .B(N2847));
INVXL inst_cellmath__60_0_I302 (.Y(N2824), .A(N2746));
NOR2XL inst_cellmath__60_0_I303 (.Y(N2779), .A(N2746), .B(N2822));
NOR2XL inst_cellmath__60_0_I304 (.Y(N2597), .A(N2746), .B(N2887));
NOR2XL inst_cellmath__60_0_I305 (.Y(N2734), .A(N2746), .B(N2637));
NOR2XL inst_cellmath__60_0_I306 (.Y(N2878), .A(N2746), .B(N2705));
NOR2XL inst_cellmath__60_0_I307 (.Y(N2694), .A(N2746), .B(N2776));
OR2XL inst_cellmath__60_0_I308 (.Y(N2711), .A(N2746), .B(N2847));
INVXL inst_cellmath__60_0_I309 (.Y(N2712), .A(N2822));
NOR2XL inst_cellmath__60_0_I310 (.Y(N2670), .A(N2822), .B(N2887));
NOR2XL inst_cellmath__60_0_I311 (.Y(N2815), .A(N2822), .B(N2637));
NOR2XL inst_cellmath__60_0_I312 (.Y(N2630), .A(N2822), .B(N2705));
NOR2XL inst_cellmath__60_0_I313 (.Y(N2771), .A(N2822), .B(N2776));
OR2XL inst_cellmath__60_0_I314 (.Y(N2783), .A(N2822), .B(N2847));
INVXL inst_cellmath__60_0_I315 (.Y(N2790), .A(N2887));
NOR2XL inst_cellmath__60_0_I316 (.Y(N2745), .A(N2887), .B(N2637));
NOR2XL inst_cellmath__60_0_I317 (.Y(N2886), .A(N2887), .B(N2705));
NOR2XL inst_cellmath__60_0_I318 (.Y(N2704), .A(N2887), .B(N2776));
OR2XL inst_cellmath__60_0_I319 (.Y(N2852), .A(N2887), .B(N2847));
INVXL inst_cellmath__60_0_I320 (.Y(N2722), .A(N2637));
NOR2XL inst_cellmath__60_0_I321 (.Y(N2681), .A(N2637), .B(N2705));
NOR2XL inst_cellmath__60_0_I322 (.Y(N2830), .A(N2637), .B(N2776));
OR2XL inst_cellmath__60_0_I323 (.Y(N2600), .A(N2637), .B(N2847));
INVXL inst_cellmath__60_0_I324 (.Y(N2842), .A(N2705));
NOR2XL inst_cellmath__60_0_I325 (.Y(N2800), .A(N2705), .B(N2776));
OR2XL inst_cellmath__60_0_I326 (.Y(N2668), .A(N2705), .B(N2847));
INVXL inst_cellmath__60_0_I327 (.Y(N2820), .A(N2776));
ADDHX1 inst_cellmath__60_0_I328 (.CO(N2813), .S(N2738), .A(N2807), .B(N2675));
ADDHX1 inst_cellmath__60_0_I329 (.CO(N2626), .S(N2881), .A(N2629), .B(N2821));
ADDHX1 inst_cellmath__60_0_I330 (.CO(N2769), .S(N2697), .A(N2616), .B(N2636));
ADDFX1 inst_cellmath__60_0_I331 (.CO(N2589), .S(N2841), .A(N2770), .B(N2762), .CI(N2626));
ADDHX1 inst_cellmath__60_0_I332 (.CO(N2726), .S(N2656), .A(N2585), .B(N2778));
ADDFX1 inst_cellmath__60_0_I333 (.CO(N2865), .S(N2799), .A(N2769), .B(N2590), .CI(N2656));
ADDHX1 inst_cellmath__60_0_I334 (.CO(N2684), .S(N2615), .A(N2609), .B(N2595));
ADDFX1 inst_cellmath__60_0_I335 (.CO(N2832), .S(N2754), .A(N2727), .B(N2578), .CI(N2721));
ADDFX1 inst_cellmath__60_0_I336 (.CO(N2645), .S(N2577), .A(N2615), .B(N2726), .CI(N2754));
ADDHX1 inst_cellmath__60_0_I337 (.CO(N2788), .S(N2714), .A(N2715), .B(N2732));
ADDFX1 inst_cellmath__60_0_I338 (.CO(N2605), .S(N2854), .A(N2867), .B(N2861), .CI(N2684));
ADDFX1 inst_cellmath__60_0_I339 (.CO(N2742), .S(N2672), .A(N2832), .B(N2714), .CI(N2854));
ADDHX1 inst_cellmath__60_0_I340 (.CO(N2885), .S(N2818), .A(N2787), .B(N2877));
ADDFX1 inst_cellmath__60_0_I341 (.CO(N2702), .S(N2633), .A(N2685), .B(N2891), .CI(N2680));
ADDFX1 inst_cellmath__60_0_I342 (.CO(N2845), .S(N2774), .A(N2788), .B(N2855), .CI(N2818));
ADDFX1 inst_cellmath__60_0_I343 (.CO(N2660), .S(N2592), .A(N2633), .B(N2605), .CI(N2774));
ADDHX1 inst_cellmath__60_0_I344 (.CO(N2805), .S(N2730), .A(N2709), .B(N2691));
ADDFX1 inst_cellmath__60_0_I345 (.CO(N2619), .S(N2871), .A(N2833), .B(N2673), .CI(N2829));
ADDFX1 inst_cellmath__60_0_I346 (.CO(N2759), .S(N2688), .A(N2730), .B(N2885), .CI(N2702));
ADDFX1 inst_cellmath__60_0_I347 (.CO(N2583), .S(N2836), .A(N2845), .B(N2871), .CI(N2688));
ADDHX1 inst_cellmath__60_0_I348 (.CO(N2719), .S(N2650), .A(N2824), .B(N2838));
ADDFX1 inst_cellmath__60_0_I349 (.CO(N2858), .S(N2793), .A(N2647), .B(N2741), .CI(N2643));
ADDFX1 inst_cellmath__60_0_I350 (.CO(N2677), .S(N2608), .A(N2819), .B(N2850), .CI(N2805));
ADDFX1 inst_cellmath__60_0_I351 (.CO(N2826), .S(N2749), .A(N2619), .B(N2650), .CI(N2793));
ADDFX1 inst_cellmath__60_0_I352 (.CO(N2639), .S(N2890), .A(N2759), .B(N2608), .CI(N2749));
XNOR2X1 inst_cellmath__60_0_I353 (.Y(N2708), .A(N2884), .B(N2789));
OR2XL inst_cellmath__60_0_I354 (.Y(N2781), .A(N2884), .B(N2789));
ADDFX1 inst_cellmath__60_0_I355 (.CO(N2735), .S(N2665), .A(N2784), .B(N2666), .CI(N2635));
ADDFX1 inst_cellmath__60_0_I356 (.CO(N2879), .S(N2809), .A(N2719), .B(N2611), .CI(N2708));
ADDFX1 inst_cellmath__60_0_I357 (.CO(N2695), .S(N2623), .A(N2677), .B(N2858), .CI(N2665));
ADDFX1 inst_cellmath__60_0_I358 (.CO(N2840), .S(N2766), .A(N2826), .B(N2809), .CI(N2623));
ADDFX1 inst_cellmath__60_0_I359 (.CO(N2655), .S(N2587), .A(N2779), .B(N2712), .CI(N2602));
ADDFX1 inst_cellmath__60_0_I360 (.CO(N2797), .S(N2724), .A(N2775), .B(N2701), .CI(N2811));
ADDFX1 inst_cellmath__60_0_I361 (.CO(N2614), .S(N2864), .A(N2781), .B(N2679), .CI(N2735));
ADDFX1 inst_cellmath__60_0_I362 (.CO(N2753), .S(N2683), .A(N2724), .B(N2587), .CI(N2879));
ADDFX1 inst_cellmath__60_0_I363 (.CO(N2895), .S(N2831), .A(N2695), .B(N2864), .CI(N2683));
ADDFX1 inst_cellmath__60_0_I364 (.CO(N2713), .S(N2644), .A(N2593), .B(N2597), .CI(N2624));
ADDFX1 inst_cellmath__60_0_I365 (.CO(N2853), .S(N2786), .A(N2752), .B(N2844), .CI(N2655));
ADDFX1 inst_cellmath__60_0_I366 (.CO(N2671), .S(N2604), .A(N2644), .B(N2797), .CI(N2614));
ADDFX1 inst_cellmath__60_0_I367 (.CO(N2816), .S(N2740), .A(N2753), .B(N2786), .CI(N2604));
ADDFX1 inst_cellmath__60_0_I368 (.CO(N2632), .S(N2883), .A(N2670), .B(N2790), .CI(N2767));
ADDFX1 inst_cellmath__60_0_I369 (.CO(N2773), .S(N2699), .A(N2659), .B(N2734), .CI(N2828));
ADDFX1 inst_cellmath__60_0_I370 (.CO(N2591), .S(N2843), .A(N2883), .B(N2713), .CI(N2699));
ADDFX1 inst_cellmath__60_0_I371 (.CO(N2729), .S(N2658), .A(N2671), .B(N2853), .CI(N2843));
ADDFX1 inst_cellmath__60_0_I372 (.CO(N2869), .S(N2801), .A(N2803), .B(N2815), .CI(N2878));
ADDFX1 inst_cellmath__60_0_I373 (.CO(N2686), .S(N2617), .A(N2632), .B(N2893), .CI(N2773));
ADDFX1 inst_cellmath__60_0_I374 (.CO(N2834), .S(N2757), .A(N2591), .B(N2801), .CI(N2617));
ADDFX1 inst_cellmath__60_0_I375 (.CO(N2649), .S(N2581), .A(N2745), .B(N2722), .CI(N2694));
ADDFX1 inst_cellmath__60_0_I376 (.CO(N2791), .S(N2717), .A(N2642), .B(N2630), .CI(N2869));
ADDFX1 inst_cellmath__60_0_I377 (.CO(N2606), .S(N2857), .A(N2686), .B(N2581), .CI(N2717));
ADDFX1 inst_cellmath__60_0_I378 (.CO(N2747), .S(N2674), .A(N2771), .B(N2886), .CI(N2711));
ADDFX1 inst_cellmath__60_0_I379 (.CO(N2888), .S(N2823), .A(N2674), .B(N2649), .CI(N2791));
ADDFX1 inst_cellmath__60_0_I380 (.CO(N2706), .S(N2638), .A(N2681), .B(N2842), .CI(N2704));
ADDFX1 inst_cellmath__60_0_I381 (.CO(N2848), .S(N2777), .A(N2747), .B(N2783), .CI(N2638));
ADDFX1 inst_cellmath__60_0_I382 (.CO(N2663), .S(N2596), .A(N2852), .B(N2830), .CI(N2706));
ADDFX1 inst_cellmath__60_0_I383 (.CO(N2808), .S(N2733), .A(N2800), .B(N2820), .CI(N2600));
AND2XL inst_cellmath__60_0_I386 (.Y(N2763), .A(N2814), .B(N2738));
NOR2XL inst_cellmath__60_0_I387 (.Y(N2839), .A(N2813), .B(N2881));
NAND2XL inst_cellmath__60_0_I388 (.Y(N2586), .A(N2813), .B(N2881));
AND2XL inst_cellmath__60_0_I390 (.Y(N2723), .A(N2697), .B(N2841));
NOR2XL inst_cellmath__60_0_I391 (.Y(N2796), .A(N2589), .B(N2799));
NAND2XL inst_cellmath__60_0_I392 (.Y(N2862), .A(N2589), .B(N2799));
AND2XL inst_cellmath__60_0_I394 (.Y(N2682), .A(N2865), .B(N2577));
NOR3XL inst_cellmath__60_0_I4935 (.Y(N2894), .A(N2631), .B(N2875), .C(N2698));
OAI22XL inst_cellmath__60_0_I4906 (.Y(N2628), .A0(N2763), .A1(N2894), .B0(N2814), .B1(N2738));
AOI21XL inst_cellmath__60_0_I399 (.Y(N2868), .A0(N2586), .A1(N2628), .B0(N2839));
OAI22XL inst_cellmath__60_0_I4907 (.Y(N2744), .A0(N2723), .A1(N2868), .B0(N2697), .B1(N2841));
AOI21XL inst_cellmath__60_0_I403 (.Y(N2621), .A0(N2862), .A1(N2744), .B0(N2796));
OAI22XL inst_cellmath__60_0_I4908 (.Y(N2846), .A0(N2682), .A1(N2621), .B0(N2865), .B1(N2577));
NOR2XL inst_cellmath__60_0_I419 (.Y(N2661), .A(N2645), .B(N2672));
XOR2XL inst_cellmath__60_0_I420 (.Y(N2731), .A(N2645), .B(N2672));
NOR2XL inst_cellmath__60_0_I421 (.Y(N2806), .A(N2742), .B(N2592));
XOR2XL inst_cellmath__60_0_I422 (.Y(N2874), .A(N2742), .B(N2592));
NOR2XL inst_cellmath__60_0_I423 (.Y(N2620), .A(N2660), .B(N2836));
XOR2XL inst_cellmath__60_0_I424 (.Y(N2689), .A(N2660), .B(N2836));
NOR2XL inst_cellmath__60_0_I425 (.Y(N2761), .A(N2583), .B(N2890));
XOR2XL inst_cellmath__60_0_I426 (.Y(N2837), .A(N2583), .B(N2890));
NOR2XL inst_cellmath__60_0_I427 (.Y(N2584), .A(N2639), .B(N2766));
XOR2XL inst_cellmath__60_0_I428 (.Y(N2652), .A(N2639), .B(N2766));
NOR2XL inst_cellmath__60_0_I429 (.Y(N2720), .A(N2840), .B(N2831));
XOR2XL inst_cellmath__60_0_I430 (.Y(N2794), .A(N2840), .B(N2831));
NOR2XL inst_cellmath__60_0_I431 (.Y(N2860), .A(N2895), .B(N2740));
XOR2XL inst_cellmath__60_0_I432 (.Y(N2610), .A(N2895), .B(N2740));
NOR2XL inst_cellmath__60_0_I433 (.Y(N2678), .A(N2816), .B(N2658));
XOR2XL inst_cellmath__60_0_I434 (.Y(N2751), .A(N2816), .B(N2658));
NOR2XL inst_cellmath__60_0_I435 (.Y(N2827), .A(N2729), .B(N2757));
XOR2XL inst_cellmath__60_0_I436 (.Y(N2892), .A(N2729), .B(N2757));
NOR2XL inst_cellmath__60_0_I437 (.Y(N2641), .A(N2834), .B(N2857));
XOR2XL inst_cellmath__60_0_I438 (.Y(N2710), .A(N2834), .B(N2857));
NOR2XL inst_cellmath__60_0_I439 (.Y(N2782), .A(N2823), .B(N2606));
XOR2XL inst_cellmath__60_0_I440 (.Y(N2851), .A(N2823), .B(N2606));
NOR2XL inst_cellmath__60_0_I441 (.Y(N2599), .A(N2888), .B(N2777));
XOR2XL inst_cellmath__60_0_I442 (.Y(N2667), .A(N2888), .B(N2777));
NOR2XL inst_cellmath__60_0_I443 (.Y(N2737), .A(N2596), .B(N2848));
XOR2XL inst_cellmath__60_0_I444 (.Y(N2812), .A(N2596), .B(N2848));
NOR2XL inst_cellmath__60_0_I445 (.Y(N2880), .A(N2733), .B(N2663));
XOR2XL inst_cellmath__60_0_I446 (.Y(N2625), .A(N2733), .B(N2663));
NOR2XL inst_cellmath__60_0_I447 (.Y(N2696), .A(N2668), .B(N2808));
XOR2XL inst_cellmath__60_0_I448 (.Y(N2768), .A(N2668), .B(N2808));
NAND2BXL inst_cellmath__60_0_I449 (.Y(N2588), .AN(N2847), .B(N2776));
AO21XL inst_cellmath__60_0_I450 (.Y(N2798), .A0(N2731), .A1(N2846), .B0(N2661));
AO21XL inst_cellmath__60_0_I451 (.Y(N2576), .A0(N2874), .A1(N2798), .B0(N2806));
AO21XL inst_cellmath__60_0_I452 (.Y(N2817), .A0(N2689), .A1(N2576), .B0(N2620));
AO21XL inst_cellmath__60_0_I453 (.Y(N2870), .A0(N2837), .A1(N2817), .B0(N2761));
AO21XL inst_cellmath__60_0_I454 (.Y(N2748), .A0(N2652), .A1(N2870), .B0(N2584));
AO21XL inst_cellmath__60_0_I455 (.Y(N2765), .A0(N2794), .A1(N2748), .B0(N2720));
AO21XL inst_cellmath__60_0_I456 (.Y(N2603), .A0(N2610), .A1(N2765), .B0(N2860));
AO21XL inst_cellmath__60_0_I457 (.Y(N2580), .A0(N2751), .A1(N2603), .B0(N2678));
AO21XL inst_cellmath__60_0_I458 (.Y(N2690), .A0(N2892), .A1(N2580), .B0(N2827));
AO21XL inst_cellmath__60_0_I459 (.Y(N2627), .A0(N2710), .A1(N2690), .B0(N2641));
AO21XL inst_cellmath__60_0_I460 (.Y(N2703), .A0(N2851), .A1(N2627), .B0(N2782));
AO21XL inst_cellmath__60_0_I461 (.Y(N2601), .A0(N2667), .A1(N2703), .B0(N2599));
AO21XL inst_cellmath__60_0_I462 (.Y(N2634), .A0(N2812), .A1(N2601), .B0(N2737));
AO21XL inst_cellmath__60_0_I463 (.Y(N2810), .A0(N2625), .A1(N2634), .B0(N2880));
AO21XL inst_cellmath__60_0_I464 (.Y(N2802), .A0(N2768), .A1(N2810), .B0(N2696));
INVXL cynw_cm_float_rcp_I481 (.Y(N3344), .A(a_man[16]));
INVXL cynw_cm_float_rcp_I482 (.Y(N3721), .A(a_man[17]));
AOI22X1 cynw_cm_float_rcp_I483 (.Y(N3480), .A0(N3344), .A1(a_man[17]), .B0(N3721), .B1(a_man[16]));
NAND2X1 cynw_cm_float_rcp_I484 (.Y(N3867), .A(N3721), .B(N3344));
NAND2X1 cynw_cm_float_rcp_I485 (.Y(N3342), .A(N3721), .B(a_man[16]));
NOR2X1 cynw_cm_float_rcp_I486 (.Y(N3750), .A(N3721), .B(N3344));
NAND2X1 cynw_cm_float_rcp_I487 (.Y(N3220), .A(a_man[16]), .B(a_man[17]));
NOR2X1 cynw_cm_float_rcp_I488 (.Y(N3634), .A(N3721), .B(a_man[16]));
NOR2XL cynw_cm_float_rcp_I489 (.Y(N4034), .A(a_man[17]), .B(a_man[16]));
NOR2XL cynw_cm_float_rcp_I490 (.Y(N3515), .A(a_man[17]), .B(N3344));
INVX3 cynw_cm_float_rcp_I491 (.Y(N3639), .A(a_man[18]));
AOI22XL cynw_cm_float_rcp_I492 (.Y(N3921), .A0(N3639), .A1(N3867), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I493 (.Y(N3855), .A0(N3639), .A1(N3634), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I494 (.Y(N4056), .A0(N3639), .A1(N3220), .B0(N3867), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I495 (.Y(N3388), .A(a_man[18]), .B(N3750));
AOI22XL cynw_cm_float_rcp_I496 (.Y(N3380), .A0(N3639), .A1(N3750), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I497 (.Y(N3581), .A0(N3639), .A1(N3721), .B0(a_man[16]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I498 (.Y(N3787), .A(N3342));
AOI22XL cynw_cm_float_rcp_I499 (.Y(N3800), .A0(N3639), .A1(N3342), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I500 (.Y(N3267), .A0(N3639), .A1(a_man[17]), .B0(a_man[16]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I501 (.Y(N3486), .A(N3480));
AOI22XL cynw_cm_float_rcp_I502 (.Y(N3670), .A0(N3639), .A1(N3634), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I503 (.Y(N4089), .A0(N3639), .A1(N3721), .B0(N3750), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I504 (.Y(N4071), .A(N3639), .B(N3220));
AOI22XL cynw_cm_float_rcp_I505 (.Y(N3598), .A0(N3639), .A1(N3634), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I506 (.Y(N4001), .A0(N3639), .A1(a_man[16]), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I507 (.Y(N3560), .A0(N3639), .A1(N3220), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I508 (.Y(N3967), .A0(N3639), .A1(N4034), .B0(a_man[17]), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I509 (.Y(N3687), .A(a_man[18]), .B(N3634));
AOI22XL cynw_cm_float_rcp_I510 (.Y(N3362), .A0(N3639), .A1(a_man[16]), .B0(N3867), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I511 (.Y(N3563), .A(N3639), .B(N3750));
NOR2XL cynw_cm_float_rcp_I512 (.Y(N3440), .A(a_man[18]), .B(N3515));
AOI22XL cynw_cm_float_rcp_I514 (.Y(N3533), .A0(N3639), .A1(N3721), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I515 (.Y(N3734), .A0(N3639), .A1(N3750), .B0(N3867), .B1(a_man[18]));
NAND2X1 cynw_cm_float_rcp_I516 (.Y(N3706), .A(N3344), .B(a_man[17]));
AOI22X1 cynw_cm_float_rcp_I517 (.Y(N3463), .A0(a_man[16]), .A1(a_man[17]), .B0(N3721), .B1(N3344));
NOR2XL cynw_cm_float_rcp_I518 (.Y(N4135), .A(N3639), .B(N4034));
AOI22XL cynw_cm_float_rcp_I519 (.Y(N3612), .A0(N3639), .A1(a_man[17]), .B0(N3721), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I520 (.Y(N4013), .A(a_man[17]), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I521 (.Y(N3492), .A0(N3639), .A1(N3463), .B0(N3706), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I522 (.Y(N3484), .A(N3639), .B(N3344));
AOI22XL cynw_cm_float_rcp_I523 (.Y(N3889), .A0(N3639), .A1(N3480), .B0(N3220), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I524 (.Y(N4097), .A0(N3639), .A1(N3220), .B0(N3463), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I525 (.Y(N3367), .A0(N3639), .A1(N3750), .B0(N3463), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I526 (.Y(N3897), .A0(N3639), .A1(a_man[16]), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I527 (.Y(N3242), .A0(N3639), .A1(N3463), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I528 (.Y(N3448), .A0(N3639), .A1(N3706), .B0(N3515), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I529 (.Y(N3393), .A(N3463));
AOI22XL cynw_cm_float_rcp_I530 (.Y(N3777), .A0(N3639), .A1(N3867), .B0(N4034), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I531 (.Y(N3248), .A(a_man[18]), .B(N3867));
NAND2XL cynw_cm_float_rcp_I532 (.Y(N3664), .A(N3639), .B(N4034));
NAND2XL cynw_cm_float_rcp_I533 (.Y(N3908), .A(N3344), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I534 (.Y(N4063), .A0(N3639), .A1(a_man[17]), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I535 (.Y(N3583), .A0(N3639), .A1(N4034), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I536 (.Y(N3541), .A0(N3639), .A1(a_man[17]), .B0(N3515), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I537 (.Y(N3987), .A(N3639), .B(a_man[17]));
NAND2XL cynw_cm_float_rcp_I538 (.Y(N3461), .A(N3639), .B(a_man[16]));
AOI22XL cynw_cm_float_rcp_I539 (.Y(N3345), .A0(N3639), .A1(N3867), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I540 (.Y(N3546), .A0(N3639), .A1(a_man[17]), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I541 (.Y(N3752), .A0(N3639), .A1(N3634), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I542 (.Y(N3947), .A0(N3639), .A1(a_man[17]), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I543 (.Y(N3427), .A0(N3639), .A1(N3463), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I544 (.Y(N3636), .A0(N3639), .A1(N3750), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I545 (.Y(N3417), .A0(N3639), .A1(N3344), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I546 (.Y(N3828), .A0(N3639), .A1(N3480), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I547 (.Y(N3299), .A0(N3639), .A1(N4034), .B0(N3867), .B1(a_man[18]));
CLKINVX6 cynw_cm_float_rcp_I550 (.Y(N3712), .A(a_man[19]));
AOI22XL cynw_cm_float_rcp_I551 (.Y(N3768), .A0(N3712), .A1(N4135), .B0(N3921), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I552 (.Y(N3969), .A0(N3712), .A1(N3344), .B0(N3855), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I554 (.Y(N3238), .A0(N3712), .A1(a_man[17]), .B0(N4056), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I555 (.Y(N3445), .A0(N3712), .A1(N3612), .B0(N3388), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I556 (.Y(N3653), .A(N3712), .B(N4013));
AOI22XL cynw_cm_float_rcp_I557 (.Y(N3405), .A0(N3712), .A1(N3492), .B0(N3380), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I558 (.Y(N3617), .A0(N3712), .A1(N3484), .B0(N3581), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I559 (.Y(N3819), .A0(N3712), .A1(N3889), .B0(N3787), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I560 (.Y(N4018), .A0(N3712), .A1(N4097), .B0(N3800), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I561 (.Y(N3289), .A0(N3712), .A1(N3367), .B0(N3267), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I562 (.Y(N3498), .A0(N3712), .A1(N3897), .B0(N3486), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I563 (.Y(N3702), .A0(N3712), .A1(N3267), .B0(N3670), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I564 (.Y(N3904), .A0(N3712), .A1(N3897), .B0(N4089), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I565 (.Y(N4111), .A0(N3712), .A1(N3242), .B0(N4071), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I566 (.Y(N3378), .A0(N3712), .A1(N3448), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I567 (.Y(N3577), .A0(N3712), .A1(N3393), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I568 (.Y(N3781), .A0(N3712), .A1(N3777), .B0(a_man[18]), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I569 (.Y(N3982), .A(a_man[19]), .B(N3248));
NOR2XL cynw_cm_float_rcp_I570 (.Y(N3709), .A(a_man[19]), .B(N3664));
AOI22XL cynw_cm_float_rcp_I571 (.Y(N3834), .A0(N3712), .A1(N2381), .B0(N3598), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I572 (.Y(N4032), .A0(N3712), .A1(N3908), .B0(N3800), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I573 (.Y(N3306), .A0(N3712), .A1(N4063), .B0(N4001), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I574 (.Y(N3513), .A0(N3712), .A1(N3583), .B0(N3560), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I575 (.Y(N3716), .A0(N3712), .A1(N3541), .B0(N3967), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I576 (.Y(N3920), .A0(N3712), .A1(N3987), .B0(N3687), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I577 (.Y(N4122), .A0(N3712), .A1(N3461), .B0(N3362), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I578 (.Y(N3386), .A0(N3712), .A1(N3967), .B0(N3563), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I579 (.Y(N3592), .A0(N3712), .A1(N4063), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I580 (.Y(N3798), .A0(N3712), .A1(N3345), .B0(N2381), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I581 (.Y(N3995), .A0(N3712), .A1(N3546), .B0(N3486), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I582 (.Y(N3265), .A0(N3712), .A1(N3752), .B0(N3533), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I583 (.Y(N3474), .A0(N3712), .A1(N3541), .B0(N3734), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I584 (.Y(N3682), .A0(N3712), .A1(N3947), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I585 (.Y(N3881), .A0(N3712), .A1(N3427), .B0(N2381), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I586 (.Y(N4087), .A(N3712), .B(N3636));
NOR2XL cynw_cm_float_rcp_I587 (.Y(N3558), .A(a_man[19]), .B(N4135));
AOI22XL cynw_cm_float_rcp_I588 (.Y(N3234), .A0(N3712), .A1(N3417), .B0(N3344), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I589 (.Y(N3439), .A0(N3712), .A1(N3828), .B0(N3721), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I590 (.Y(N3648), .A0(N3712), .A1(N3299), .B0(N3639), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I591 (.Y(N3848), .A(N3712), .B(N3664));
NAND2XL cynw_cm_float_rcp_I592 (.Y(N3324), .A(N3712), .B(N3248));
NOR2XL cynw_cm_float_rcp_I593 (.Y(N4118), .A(N3639), .B(N3721));
AOI22XL cynw_cm_float_rcp_I594 (.Y(N3588), .A0(N3639), .A1(N3867), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I595 (.Y(N3990), .A0(N3639), .A1(N3634), .B0(N3515), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I596 (.Y(N3755), .A0(N3639), .A1(N3220), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I597 (.Y(N3955), .A0(N3639), .A1(N4034), .B0(a_man[16]), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I598 (.Y(N4039), .A(a_man[18]), .B(N4034));
AOI22XL cynw_cm_float_rcp_I599 (.Y(N3467), .A0(N3639), .A1(a_man[16]), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I600 (.Y(N3874), .A0(N3639), .A1(N3463), .B0(N3721), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I601 (.Y(N3350), .A0(N3639), .A1(N3706), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I602 (.Y(N3759), .A0(N3639), .A1(N3480), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I603 (.Y(N3227), .A0(N3639), .A1(N3750), .B0(N3721), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I604 (.Y(N3641), .A(N3639), .B(N3220));
AOI22XL cynw_cm_float_rcp_I605 (.Y(N3771), .A0(N3639), .A1(a_man[16]), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I606 (.Y(N3971), .A0(N3639), .A1(N3515), .B0(N3220), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I607 (.Y(N3240), .A(N3639), .B(N3867));
NOR2XL cynw_cm_float_rcp_I608 (.Y(N3854), .A(a_man[18]), .B(N3220));
AOI22XL cynw_cm_float_rcp_I609 (.Y(N4044), .A0(N3639), .A1(N3463), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I610 (.Y(N3938), .A0(N3639), .A1(N3706), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I611 (.Y(N3524), .A0(N3639), .A1(N3342), .B0(N3463), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I612 (.Y(N3703), .A0(N3639), .A1(N3706), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I613 (.Y(N3931), .A0(N3639), .A1(N3750), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I614 (.Y(N3397), .A0(N3639), .A1(N3515), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I615 (.Y(N3809), .A0(N3639), .A1(a_man[16]), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I616 (.Y(N3785), .A0(N3639), .A1(N3721), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I617 (.Y(N3277), .A0(N3639), .A1(N3721), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I618 (.Y(N3349), .A0(N3639), .A1(N3344), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I619 (.Y(N4132), .A0(N3639), .A1(N3750), .B0(N3220), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I620 (.Y(N3691), .A0(N3639), .A1(N3867), .B0(N3721), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I621 (.Y(N3606), .A(N3867));
AOI22XL cynw_cm_float_rcp_I622 (.Y(N3808), .A0(N3639), .A1(N3515), .B0(N3750), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I623 (.Y(N4006), .A(N4034), .B(a_man[18]));
NAND2XL cynw_cm_float_rcp_I624 (.Y(N4100), .A(N3639), .B(N3706));
AOI22XL cynw_cm_float_rcp_I625 (.Y(N3891), .A0(N3639), .A1(N3721), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I626 (.Y(N4099), .A0(N3639), .A1(N3721), .B0(N3463), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I627 (.Y(N3568), .A0(N3639), .A1(N3634), .B0(N3463), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I628 (.Y(N3974), .A0(N3639), .A1(N3342), .B0(N3515), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I629 (.Y(N3450), .A(N3867), .B(a_man[18]));
NOR2XL cynw_cm_float_rcp_I630 (.Y(N3622), .A(N3639), .B(a_man[16]));
NAND2XL cynw_cm_float_rcp_I631 (.Y(N3503), .A(N3639), .B(N3342));
AOI22XL cynw_cm_float_rcp_I632 (.Y(N3585), .A0(N3639), .A1(a_man[16]), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I633 (.Y(N3792), .A0(N3639), .A1(N3750), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I634 (.Y(N3464), .A0(N3639), .A1(N3706), .B0(N3220), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I635 (.Y(N3872), .A(N3639), .B(N3515));
AOI22XL cynw_cm_float_rcp_I636 (.Y(N3858), .A0(N3639), .A1(N3706), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I637 (.Y(N3927), .A0(N3639), .A1(a_man[17]), .B0(N3463), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I638 (.Y(N3333), .A(N3639), .B(N3750));
NAND2XL cynw_cm_float_rcp_I639 (.Y(N3241), .A(N3712), .B(N3987));
AOI22XL cynw_cm_float_rcp_I640 (.Y(N3656), .A0(N3712), .A1(N3349), .B0(N3344), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I641 (.Y(N3856), .A0(N3712), .A1(N3874), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I642 (.Y(N4057), .A0(N3712), .A1(N3227), .B0(N3612), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I643 (.Y(N3331), .A0(N3712), .A1(N4013), .B0(N4118), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I644 (.Y(N3536), .A(N3712), .B(N4013));
AOI22XL cynw_cm_float_rcp_I645 (.Y(N3292), .A0(N3712), .A1(N4132), .B0(N3588), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I646 (.Y(N3501), .A0(N3712), .A1(N3691), .B0(N3990), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I647 (.Y(N3705), .A0(N3712), .A1(N3606), .B0(N3755), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I648 (.Y(N3907), .A0(N3712), .A1(N3808), .B0(N3955), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I649 (.Y(N4114), .A0(N3712), .A1(N4006), .B0(N3560), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I650 (.Y(N3381), .A0(N3712), .A1(N4100), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I651 (.Y(N3582), .A0(N3712), .A1(N3891), .B0(N4039), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I652 (.Y(N3788), .A0(N3712), .A1(N4099), .B0(N3467), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I653 (.Y(N3986), .A0(N3712), .A1(N3427), .B0(N3874), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I654 (.Y(N3256), .A0(N3712), .A1(N3568), .B0(N3350), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I655 (.Y(N3460), .A0(N3712), .A1(N3974), .B0(N3759), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I656 (.Y(N3671), .A0(N3712), .A1(N3277), .B0(N3227), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I657 (.Y(N3870), .A0(N3712), .A1(N3450), .B0(N3641), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I658 (.Y(N3741), .A(N3712), .B(N3450));
AOI22XL cynw_cm_float_rcp_I659 (.Y(N3312), .A0(N3712), .A1(N3622), .B0(N3771), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I660 (.Y(N3519), .A0(N3712), .A1(N4044), .B0(N3971), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I661 (.Y(N3720), .A0(N3712), .A1(N3503), .B0(N3240), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I662 (.Y(N3925), .A0(N3712), .A1(N4135), .B0(N3854), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I663 (.Y(N4128), .A0(N3712), .A1(N3585), .B0(N3800), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I664 (.Y(N3391), .A0(N3712), .A1(N3792), .B0(N4044), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I665 (.Y(N3600), .A0(N3712), .A1(N3345), .B0(N3938), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I666 (.Y(N3805), .A0(N3712), .A1(N3588), .B0(N3560), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I667 (.Y(N4002), .A0(N3712), .A1(N3464), .B0(N4089), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I668 (.Y(N3272), .A0(N3712), .A1(N3809), .B0(N3524), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I669 (.Y(N3479), .A0(N3712), .A1(N3872), .B0(N3524), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I670 (.Y(N3688), .A(N3712), .B(N3858));
AOI22XL cynw_cm_float_rcp_I671 (.Y(N4093), .A0(N3712), .A1(N3921), .B0(N3955), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I672 (.Y(N3363), .A0(N3712), .A1(a_man[17]), .B0(N3703), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I673 (.Y(N3564), .A0(N3712), .A1(N2381), .B0(N3931), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I674 (.Y(N3767), .A0(N3712), .A1(N3344), .B0(N3397), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I675 (.Y(N3968), .A0(N3712), .A1(N3721), .B0(N4063), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I676 (.Y(N3236), .A0(N3712), .A1(N3467), .B0(N3809), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I677 (.Y(N3443), .A0(N3712), .A1(N3927), .B0(N3785), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I678 (.Y(N3651), .A0(N3712), .A1(N3333), .B0(N3277), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I679 (.Y(N3852), .A0(N3712), .A1(a_man[18]), .B0(N2381), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I680 (.Y(N4052), .A(a_man[19]), .B(a_man[18]));
NAND2XL cynw_cm_float_rcp_I681 (.Y(N3735), .A(N3712), .B(N3639));
INVX3 cynw_cm_float_rcp_I682 (.Y(N3409), .A(a_man[20]));
AOI22XL cynw_cm_float_rcp_I683 (.Y(N3818), .A0(N3409), .A1(N3241), .B0(N3768), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I684 (.Y(N4017), .A0(N3409), .A1(N3656), .B0(N3969), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I685 (.Y(N3288), .A0(N3409), .A1(N3856), .B0(N3238), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I686 (.Y(N3497), .A0(N3409), .A1(N4057), .B0(N3445), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I687 (.Y(N3700), .A0(N3409), .A1(N3331), .B0(N3653), .B1(a_man[20]));
NOR2XL cynw_cm_float_rcp_I688 (.Y(N3902), .A(a_man[20]), .B(N3536));
AOI22XL cynw_cm_float_rcp_I689 (.Y(N4067), .A0(N3409), .A1(N3292), .B0(N3405), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I690 (.Y(N3339), .A0(N3409), .A1(N3501), .B0(N3617), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I691 (.Y(N3544), .A0(N3409), .A1(N3705), .B0(N3819), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I692 (.Y(N3747), .A0(N3409), .A1(N3907), .B0(N4018), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I693 (.Y(N3950), .A0(N3409), .A1(N4114), .B0(N3289), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I694 (.Y(N3218), .A0(N3409), .A1(N3381), .B0(N3498), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I695 (.Y(N3423), .A0(N3409), .A1(N3582), .B0(N3702), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I696 (.Y(N3632), .A0(N3409), .A1(N3788), .B0(N3904), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I697 (.Y(N3833), .A0(N3409), .A1(N3986), .B0(N4111), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I698 (.Y(N4031), .A0(N3409), .A1(N3256), .B0(N3378), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I699 (.Y(N3304), .A0(N3409), .A1(N3460), .B0(N3577), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I700 (.Y(N3511), .A0(N3409), .A1(N3671), .B0(N3781), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I701 (.Y(N3714), .A0(N3409), .A1(N3870), .B0(N3982), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I702 (.Y(N3918), .A0(N3409), .A1(N3741), .B0(N3709), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I703 (.Y(N4120), .A(N3409), .B(N3558));
AOI22XL cynw_cm_float_rcp_I704 (.Y(N3472), .A0(N3409), .A1(N3312), .B0(N3834), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I705 (.Y(N3680), .A0(N3409), .A1(N3519), .B0(N4032), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I706 (.Y(N3879), .A0(N3409), .A1(N3720), .B0(N3306), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I707 (.Y(N4085), .A0(N3409), .A1(N3925), .B0(N3513), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I708 (.Y(N3355), .A0(N3409), .A1(N4128), .B0(N3716), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I709 (.Y(N3556), .A0(N3409), .A1(N3391), .B0(N3920), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I710 (.Y(N3764), .A0(N3409), .A1(N3600), .B0(N4122), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I711 (.Y(N3965), .A0(N3409), .A1(N3805), .B0(N3386), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I712 (.Y(N3232), .A0(N3409), .A1(N4002), .B0(N3592), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I713 (.Y(N3437), .A0(N3409), .A1(N3272), .B0(N3798), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I714 (.Y(N3646), .A0(N3409), .A1(N3479), .B0(N3995), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I715 (.Y(N3845), .A0(N3409), .A1(N3688), .B0(N3265), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I716 (.Y(N4049), .A0(N3409), .A1(N4093), .B0(N3474), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I717 (.Y(N3323), .A0(N3409), .A1(N3363), .B0(N3682), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I718 (.Y(N3530), .A0(N3409), .A1(N3564), .B0(N3881), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I719 (.Y(N3730), .A0(N3409), .A1(N3767), .B0(N4087), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I720 (.Y(N3934), .A0(N3409), .A1(N3968), .B0(N3558), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I721 (.Y(N4134), .A0(N3409), .A1(N3236), .B0(N3234), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I722 (.Y(N3399), .A0(N3409), .A1(N3443), .B0(N3439), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I723 (.Y(N3610), .A0(N3409), .A1(N3651), .B0(N3648), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I724 (.Y(N3812), .A0(N3409), .A1(N3852), .B0(N3848), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I725 (.Y(N4010), .A0(N3409), .A1(N4052), .B0(N3324), .B1(a_man[20]));
NOR2XL cynw_cm_float_rcp_I726 (.Y(N3281), .A(a_man[20]), .B(N3735));
AOI22XL cynw_cm_float_rcp_I727 (.Y(N3210), .A0(N3639), .A1(N3515), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I728 (.Y(N3790), .A0(N3639), .A1(N3706), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I729 (.Y(N3637), .A0(N3639), .A1(N3750), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I730 (.Y(N3623), .A0(N3639), .A1(N3706), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I731 (.Y(N3313), .A0(N3639), .A1(N3344), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I732 (.Y(N3520), .A0(N3639), .A1(N3750), .B0(N3706), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I733 (.Y(N3722), .A(N3639), .B(N3463));
AOI22XL cynw_cm_float_rcp_I734 (.Y(N3392), .A0(N3639), .A1(N3344), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I735 (.Y(N4023), .A0(N3639), .A1(N3463), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I736 (.Y(N3504), .A0(N3639), .A1(N3342), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I737 (.Y(N3911), .A0(N3639), .A1(a_man[17]), .B0(N3220), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I738 (.Y(N3382), .A(N3639), .B(N3721));
NOR2XL cynw_cm_float_rcp_I739 (.Y(N3737), .A(N3639), .B(N3515));
AOI22XL cynw_cm_float_rcp_I740 (.Y(N4019), .A0(N3639), .A1(N3706), .B0(N3721), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I741 (.Y(N3793), .A0(N3639), .A1(a_man[17]), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I742 (.Y(N3499), .A0(N3639), .A1(N3463), .B0(N3220), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I743 (.Y(N3579), .A0(N3639), .A1(N3706), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I744 (.Y(N3783), .A0(N3639), .A1(a_man[16]), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I745 (.Y(N3983), .A0(N3639), .A1(N3706), .B0(N4034), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I746 (.Y(N3253), .A(N3634));
AOI22XL cynw_cm_float_rcp_I747 (.Y(N3258), .A0(N3639), .A1(a_man[16]), .B0(N3463), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I748 (.Y(N3674), .A0(N3639), .A1(N3480), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I749 (.Y(N3806), .A0(N3639), .A1(N3480), .B0(N3515), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I750 (.Y(N4077), .A0(N3639), .A1(N3480), .B0(N3721), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I751 (.Y(N3487), .A0(N3639), .A1(N3344), .B0(N3634), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I752 (.Y(N3823), .A(N3639), .B(N3463));
NAND2XL cynw_cm_float_rcp_I753 (.Y(N3296), .A(N3706), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I754 (.Y(N3910), .A0(N3639), .A1(N4034), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I755 (.Y(N3584), .A0(N3639), .A1(N4034), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I756 (.Y(N3791), .A0(N3639), .A1(N3463), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I757 (.Y(N3988), .A0(N3639), .A1(N3721), .B0(N3634), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I758 (.Y(N4076), .A(N3220));
NOR2XL cynw_cm_float_rcp_I759 (.Y(N3548), .A(N3639), .B(a_man[17]));
AOI22XL cynw_cm_float_rcp_I760 (.Y(N3956), .A0(N3639), .A1(N3344), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I761 (.Y(N4040), .A0(N3639), .A1(N3721), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I762 (.Y(N3429), .A0(N3639), .A1(a_man[16]), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I763 (.Y(N3887), .A0(N3712), .A1(N3504), .B0(N3210), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I764 (.Y(N4095), .A0(N3712), .A1(N4099), .B0(N3492), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I765 (.Y(N3365), .A0(N3712), .A1(N3809), .B0(N3790), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I766 (.Y(N3566), .A0(N3712), .A1(N3793), .B0(N3277), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I767 (.Y(N3739), .A0(N3712), .A1(N3299), .B0(N3637), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I768 (.Y(N3940), .A0(N3712), .A1(N3734), .B0(N3858), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I769 (.Y(N3206), .A0(N3712), .A1(N3806), .B0(N3623), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I770 (.Y(N3407), .A0(N3712), .A1(N4077), .B0(N3313), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I771 (.Y(N3619), .A(N3712), .B(N3520));
AOI22XL cynw_cm_float_rcp_I772 (.Y(N3290), .A0(N3712), .A1(N3487), .B0(N3722), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I773 (.Y(N3500), .A0(N3712), .A1(N4089), .B0(N3392), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I774 (.Y(N3704), .A0(N3712), .A1(a_man[16]), .B0(N3277), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I775 (.Y(N3906), .A0(N3712), .A1(N3486), .B0(N3417), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I776 (.Y(N4113), .A0(N3712), .A1(N3777), .B0(N4023), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I777 (.Y(N3379), .A0(N3712), .A1(N3809), .B0(N3504), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I778 (.Y(N3580), .A0(N3712), .A1(N4023), .B0(N3947), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I779 (.Y(N3786), .A0(N3712), .A1(N3691), .B0(N3911), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I780 (.Y(N3985), .A0(N3712), .A1(N3248), .B0(N3382), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I781 (.Y(N3953), .A0(N3712), .A1(N3823), .B0(N4100), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I782 (.Y(N3222), .A0(N3712), .A1(N3296), .B0(N3641), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I783 (.Y(N3426), .A0(N3712), .A1(N3588), .B0(N3777), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I784 (.Y(N3635), .A0(N3712), .A1(N3910), .B0(N3737), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I785 (.Y(N3837), .A0(N3712), .A1(N3759), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I786 (.Y(N4037), .A0(N3712), .A1(N3623), .B0(N4019), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I787 (.Y(N3311), .A0(N3712), .A1(N3584), .B0(N3793), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I788 (.Y(N3518), .A0(N3712), .A1(N3791), .B0(N3499), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I789 (.Y(N3719), .A0(N3712), .A1(N3988), .B0(N3908), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I790 (.Y(N3924), .A0(N3712), .A1(N3579), .B0(N3382), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I791 (.Y(N4127), .A0(N3712), .A1(N3267), .B0(N3579), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I792 (.Y(N3390), .A0(N3712), .A1(N3382), .B0(N3783), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I793 (.Y(N3597), .A0(N3712), .A1(N4076), .B0(N3983), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I794 (.Y(N3803), .A0(N3712), .A1(N3908), .B0(N3253), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I795 (.Y(N4000), .A0(N3712), .A1(N3548), .B0(N3258), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I796 (.Y(N3271), .A0(N3712), .A1(N4013), .B0(N3828), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I797 (.Y(N3478), .A0(N3712), .A1(N3956), .B0(N3397), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I798 (.Y(N3686), .A0(N3712), .A1(N4040), .B0(N3674), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I799 (.Y(N3885), .A0(N3712), .A1(N3429), .B0(N3397), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I800 (.Y(N4092), .A0(N3712), .A1(N3277), .B0(N4063), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I801 (.Y(N3361), .A0(N3712), .A1(N2381), .B0(N3450), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I802 (.Y(N3412), .A(N3750), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I803 (.Y(N3838), .A0(N3639), .A1(N3344), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I804 (.Y(N4024), .A0(N3639), .A1(N3463), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I805 (.Y(N4078), .A0(N3639), .A1(N3750), .B0(a_man[16]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I806 (.Y(N3549), .A(N3706));
AOI22XL cynw_cm_float_rcp_I807 (.Y(N3430), .A0(N3639), .A1(N4034), .B0(N3463), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I808 (.Y(N3972), .A0(N3639), .A1(a_man[16]), .B0(N3515), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I809 (.Y(N3658), .A0(N3639), .A1(N3342), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I810 (.Y(N3207), .A0(N3639), .A1(N3721), .B0(N3220), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I811 (.Y(N3293), .A(N3639), .B(N3867));
AOI22XL cynw_cm_float_rcp_I812 (.Y(N4115), .A0(N3639), .A1(N3515), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I813 (.Y(N3528), .A0(N3639), .A1(N3515), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I814 (.Y(N3315), .A0(N3639), .A1(N3463), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I815 (.Y(N3608), .A0(N3639), .A1(N3220), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I816 (.Y(N3246), .A0(N3639), .A1(N4034), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I817 (.Y(N3825), .A0(N3639), .A1(N3634), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I818 (.Y(N3297), .A0(N3639), .A1(N3480), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I819 (.Y(N3757), .A0(N3639), .A1(N3342), .B0(a_man[17]), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I820 (.Y(N3958), .A(N3515));
NAND2XL cynw_cm_float_rcp_I821 (.Y(N3225), .A(N3342), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I822 (.Y(N4042), .A0(N3639), .A1(N4034), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I823 (.Y(N3317), .A0(N3639), .A1(N3634), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I824 (.Y(N3726), .A0(N3639), .A1(N3342), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I825 (.Y(N3929), .A0(N3639), .A1(N3750), .B0(N3480), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I826 (.Y(N3395), .A(a_man[18]), .B(N3344));
AOI22XL cynw_cm_float_rcp_I827 (.Y(N3724), .A0(N3639), .A1(N3220), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I828 (.Y(N3209), .A0(N3712), .A1(N3528), .B0(N3333), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I829 (.Y(N3410), .A0(N3712), .A1(N3382), .B0(N3412), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I830 (.Y(N3621), .A0(N3712), .A1(N3315), .B0(N3838), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I831 (.Y(N3822), .A0(N3712), .A1(N3568), .B0(N4024), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I832 (.Y(N4022), .A0(N3712), .A1(N3608), .B0(N3641), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I833 (.Y(N3295), .A0(N3712), .A1(N3388), .B0(N3641), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I834 (.Y(N3502), .A(N3641), .B(a_man[19]));
AOI22XL cynw_cm_float_rcp_I835 (.Y(N3257), .A0(N3712), .A1(N3806), .B0(N4078), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I836 (.Y(N3462), .A0(N3712), .A1(N3246), .B0(N3504), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I837 (.Y(N3673), .A0(N3712), .A1(N3737), .B0(N3549), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I838 (.Y(N3871), .A0(N3712), .A1(N3392), .B0(N3636), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I839 (.Y(N4075), .A0(N3712), .A1(N3737), .B0(N3858), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I840 (.Y(N3346), .A0(N3712), .A1(N3503), .B0(N3427), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I841 (.Y(N3547), .A0(N3712), .A1(N3546), .B0(N3430), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I842 (.Y(N3754), .A0(N3712), .A1(N3828), .B0(N3412), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I843 (.Y(N3954), .A(N3712), .B(N3825));
NOR2XL cynw_cm_float_rcp_I844 (.Y(N3428), .A(a_man[19]), .B(N3612));
AOI22XL cynw_cm_float_rcp_I845 (.Y(N4038), .A0(N3712), .A1(N3297), .B0(N3344), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I846 (.Y(N3314), .A0(N3712), .A1(N3568), .B0(N3393), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I847 (.Y(N3521), .A0(N3712), .A1(N4063), .B0(N3777), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I848 (.Y(N3723), .A0(N3712), .A1(N2381), .B0(N3664), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I849 (.Y(N3926), .A(a_man[19]), .B(N3382));
AOI22XL cynw_cm_float_rcp_I850 (.Y(N3481), .A0(N3712), .A1(N3333), .B0(N4071), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I851 (.Y(N3689), .A0(N3712), .A1(N3757), .B0(N3972), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I852 (.Y(N3886), .A0(N3712), .A1(N3958), .B0(N3639), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I853 (.Y(N4094), .A0(N3712), .A1(N3225), .B0(N3658), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I854 (.Y(N3364), .A0(N3712), .A1(N4001), .B0(N3974), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I855 (.Y(N3565), .A0(N3712), .A1(N3990), .B0(N3910), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I856 (.Y(N3770), .A0(N3712), .A1(N4042), .B0(N3783), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I857 (.Y(N3970), .A0(N3712), .A1(N3317), .B0(N3210), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I858 (.Y(N3239), .A0(N3712), .A1(N3956), .B0(N3947), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I859 (.Y(N3447), .A0(N3712), .A1(N3726), .B0(N3417), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I860 (.Y(N3654), .A0(N3712), .A1(N3929), .B0(N3207), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I861 (.Y(N3853), .A0(N3712), .A1(N3504), .B0(N3612), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I862 (.Y(N4055), .A0(N3712), .A1(N3395), .B0(N3670), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I863 (.Y(N3328), .A0(N3712), .A1(N3210), .B0(N3541), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I864 (.Y(N3535), .A0(N3712), .A1(N3296), .B0(N3759), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I865 (.Y(N3738), .A0(N3712), .A1(N3429), .B0(N3293), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I866 (.Y(N3937), .A0(N3712), .A1(N3674), .B0(N3467), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I867 (.Y(N3205), .A0(N3712), .A1(N3724), .B0(N4077), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I868 (.Y(N3406), .A0(N3712), .A1(N3956), .B0(N4115), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I869 (.Y(N3618), .A0(N3712), .A1(N4024), .B0(N3947), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I870 (.Y(N3820), .A0(N3712), .A1(N3641), .B0(N4135), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I871 (.Y(N4020), .A0(N3712), .A1(N3388), .B0(N4135), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I872 (.Y(N3784), .A0(N3409), .A1(N3209), .B0(N3887), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I873 (.Y(N3984), .A0(N3409), .A1(N3410), .B0(N4095), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I874 (.Y(N3254), .A0(N3409), .A1(N3621), .B0(N3365), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I875 (.Y(N3458), .A0(N3409), .A1(N3822), .B0(N3566), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I876 (.Y(N3668), .A0(N3409), .A1(N4022), .B0(N3852), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I877 (.Y(N3868), .A0(N3409), .A1(N3295), .B0(N3735), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I878 (.Y(N4069), .A(N3409), .B(N3502));
NOR2XL cynw_cm_float_rcp_I879 (.Y(N3796), .A(N3712), .B(N3388));
NOR2XL cynw_cm_float_rcp_I880 (.Y(N3952), .A(N3796), .B(a_man[20]));
AOI22XL cynw_cm_float_rcp_I881 (.Y(N4035), .A0(N3409), .A1(N3257), .B0(N3739), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I882 (.Y(N3309), .A0(N3409), .A1(N3462), .B0(N3940), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I883 (.Y(N3516), .A0(N3409), .A1(N3673), .B0(N3206), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I884 (.Y(N3717), .A0(N3409), .A1(N3871), .B0(N3407), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I885 (.Y(N3922), .A0(N3409), .A1(N4075), .B0(N3619), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I886 (.Y(N4125), .A0(N3409), .A1(N3346), .B0(N3290), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I887 (.Y(N3389), .A0(N3409), .A1(N3547), .B0(N3500), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I888 (.Y(N3595), .A0(N3409), .A1(N3754), .B0(N3704), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I889 (.Y(N3801), .A0(N3409), .A1(N3954), .B0(N3906), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I890 (.Y(N3998), .A0(N3409), .A1(N3428), .B0(N4113), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I891 (.Y(N3268), .A0(N3409), .A1(N4038), .B0(N3379), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I892 (.Y(N3476), .A0(N3409), .A1(N3314), .B0(N3580), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I893 (.Y(N3684), .A0(N3409), .A1(N3521), .B0(N3786), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I894 (.Y(N3883), .A0(N3409), .A1(N3723), .B0(N3985), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I895 (.Y(N4090), .A0(N3409), .A1(N3926), .B0(N3324), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I896 (.Y(N3649), .A0(N3409), .A1(N3481), .B0(N3953), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I897 (.Y(N3850), .A0(N3409), .A1(N3689), .B0(N3222), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I898 (.Y(N4050), .A0(N3409), .A1(N3886), .B0(N3426), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I899 (.Y(N3325), .A0(N3409), .A1(N4094), .B0(N3635), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I900 (.Y(N3531), .A0(N3409), .A1(N3364), .B0(N3837), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I901 (.Y(N3732), .A0(N3409), .A1(N3565), .B0(N4037), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I902 (.Y(N3935), .A0(N3409), .A1(N3770), .B0(N3311), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I903 (.Y(N3203), .A0(N3409), .A1(N3970), .B0(N3518), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I904 (.Y(N3403), .A0(N3409), .A1(N3239), .B0(N3719), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I905 (.Y(N3614), .A0(N3409), .A1(N3447), .B0(N3924), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I906 (.Y(N3816), .A0(N3409), .A1(N3654), .B0(N4127), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I907 (.Y(N4015), .A0(N3409), .A1(N3853), .B0(N3390), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I908 (.Y(N3285), .A0(N3409), .A1(N4055), .B0(N3597), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I909 (.Y(N3494), .A0(N3409), .A1(N3328), .B0(N3803), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I910 (.Y(N3697), .A0(N3409), .A1(N3535), .B0(N4000), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I911 (.Y(N3899), .A0(N3409), .A1(N3738), .B0(N3271), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I912 (.Y(N4107), .A0(N3409), .A1(N3937), .B0(N3478), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I913 (.Y(N3374), .A0(N3409), .A1(N3205), .B0(N3686), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I914 (.Y(N3574), .A0(N3409), .A1(N3406), .B0(N3885), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I915 (.Y(N3779), .A0(N3409), .A1(N3618), .B0(N4092), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I916 (.Y(N3979), .A0(N3409), .A1(N3820), .B0(N3361), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I917 (.Y(N3250), .A0(N3409), .A1(N4020), .B0(a_man[19]), .B1(a_man[20]));
OAI2BB1X1 cynw_cm_float_rcp_I918 (.Y(N3455), .A0N(N4135), .A1N(a_man[19]), .B0(N3409));
NOR2XL cynw_cm_float_rcp_I919 (.Y(N3356), .A(N3712), .B(N3450));
NOR2XL cynw_cm_float_rcp_I920 (.Y(N3864), .A(N3356), .B(a_man[20]));
INVX1 cynw_cm_float_rcp_I921 (.Y(N4112), .A(a_man[21]));
AOI22XL cynw_cm_float_rcp_I922 (.Y(N3216), .A0(N4112), .A1(N3784), .B0(N3818), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I923 (.Y(N3419), .A0(N4112), .A1(N3984), .B0(N4017), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I924 (.Y(N3629), .A0(N4112), .A1(N3254), .B0(N3288), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I925 (.Y(N3830), .A0(N4112), .A1(N3458), .B0(N3497), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I926 (.Y(N4027), .A0(N4112), .A1(N3668), .B0(N3700), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I927 (.Y(N3301), .A0(N4112), .A1(N3868), .B0(N3902), .B1(a_man[21]));
NAND2XL cynw_cm_float_rcp_I928 (.Y(N3508), .A(N4112), .B(N4069));
NOR2XL cynw_cm_float_rcp_I929 (.Y(N3915), .A(a_man[21]), .B(N4069));
NAND2XL cynw_cm_float_rcp_I930 (.Y(N3590), .A(N4112), .B(N3952));
AOI22XL cynw_cm_float_rcp_I931 (.Y(N3262), .A0(N4112), .A1(N4035), .B0(N4067), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I932 (.Y(N3469), .A0(N4112), .A1(N3309), .B0(N3339), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I933 (.Y(N3677), .A0(N4112), .A1(N3516), .B0(N3544), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I934 (.Y(N3876), .A0(N4112), .A1(N3717), .B0(N3747), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I935 (.Y(N4082), .A0(N4112), .A1(N3922), .B0(N3950), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I936 (.Y(N3352), .A0(N4112), .A1(N4125), .B0(N3218), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I937 (.Y(N3553), .A0(N4112), .A1(N3389), .B0(N3423), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I938 (.Y(N3761), .A0(N4112), .A1(N3595), .B0(N3632), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I939 (.Y(N3962), .A0(N4112), .A1(N3801), .B0(N3833), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I940 (.Y(N3229), .A0(N4112), .A1(N3998), .B0(N4031), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I941 (.Y(N3434), .A0(N4112), .A1(N3268), .B0(N3304), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I942 (.Y(N3643), .A0(N4112), .A1(N3476), .B0(N3511), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I943 (.Y(N3842), .A0(N4112), .A1(N3684), .B0(N3714), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I944 (.Y(N4046), .A0(N4112), .A1(N3883), .B0(N3918), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I945 (.Y(N3320), .A0(N4112), .A1(N4090), .B0(N4120), .B1(a_man[21]));
NOR2XL cynw_cm_float_rcp_I946 (.Y(N3846), .A(N3409), .B(N3709));
NOR2XL cynw_cm_float_rcp_I947 (.Y(N3526), .A(N3846), .B(a_man[21]));
AOI22XL cynw_cm_float_rcp_I948 (.Y(N3810), .A0(N4112), .A1(N3649), .B0(N3472), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I949 (.Y(N4007), .A0(N4112), .A1(N3850), .B0(N3680), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I950 (.Y(N3278), .A0(N4112), .A1(N4050), .B0(N3879), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I951 (.Y(N3488), .A0(N4112), .A1(N3325), .B0(N4085), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I952 (.Y(N3692), .A0(N4112), .A1(N3531), .B0(N3355), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I953 (.Y(N3892), .A0(N4112), .A1(N3732), .B0(N3556), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I954 (.Y(N4101), .A0(N4112), .A1(N3935), .B0(N3764), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I955 (.Y(N3369), .A0(N4112), .A1(N3203), .B0(N3965), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I956 (.Y(N3569), .A0(N4112), .A1(N3403), .B0(N3232), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I957 (.Y(N3774), .A0(N4112), .A1(N3614), .B0(N3437), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I958 (.Y(N3975), .A0(N4112), .A1(N3816), .B0(N3646), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I959 (.Y(N3244), .A0(N4112), .A1(N4015), .B0(N3845), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I960 (.Y(N3451), .A0(N4112), .A1(N3285), .B0(N4049), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I961 (.Y(N3660), .A0(N4112), .A1(N3494), .B0(N3323), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I962 (.Y(N3859), .A0(N4112), .A1(N3697), .B0(N3530), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I963 (.Y(N4060), .A0(N4112), .A1(N3899), .B0(N3730), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I964 (.Y(N3334), .A0(N4112), .A1(N4107), .B0(N3934), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I965 (.Y(N3538), .A0(N4112), .A1(N3374), .B0(N4134), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I966 (.Y(N3742), .A0(N4112), .A1(N3574), .B0(N3399), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I967 (.Y(N3943), .A0(N4112), .A1(N3779), .B0(N3610), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I968 (.Y(N3211), .A0(N4112), .A1(N3979), .B0(N3812), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I969 (.Y(N3413), .A0(N4112), .A1(N3250), .B0(N4010), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I970 (.Y(N3624), .A0(N4112), .A1(N3455), .B0(N3281), .B1(a_man[21]));
NAND2XL cynw_cm_float_rcp_I971 (.Y(N3824), .A(N4112), .B(N3864));
AOI22XL cynw_cm_float_rcp_I972 (.Y(N3616), .A0(N3639), .A1(N3344), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I973 (.Y(N3422), .A0(N3639), .A1(N3463), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I974 (.Y(N4030), .A0(N3639), .A1(N3634), .B0(N3721), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I975 (.Y(N3993), .A0(N3639), .A1(N3867), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I976 (.Y(N3941), .A0(N3639), .A1(N3706), .B0(N3463), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I977 (.Y(N3672), .A(N3721), .B(a_man[18]));
NOR2XL cynw_cm_float_rcp_I978 (.Y(N4074), .A(N3639), .B(N3344));
NAND2XL cynw_cm_float_rcp_I979 (.Y(N3753), .A(N3463), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I980 (.Y(N3769), .A0(N3639), .A1(N3867), .B0(N3220), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I981 (.Y(N3446), .A0(N3639), .A1(N3220), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I982 (.Y(N4054), .A0(N3639), .A1(a_man[17]), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I983 (.Y(N3749), .A0(N3712), .A1(N3382), .B0(N4115), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I984 (.Y(N3951), .A0(N3712), .A1(N3315), .B0(N3938), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I985 (.Y(N3219), .A0(N3712), .A1(N3921), .B0(N3492), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I986 (.Y(N3424), .A0(N3712), .A1(N3941), .B0(N3790), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I987 (.Y(N3633), .A0(N3712), .A1(N3207), .B0(N4063), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I988 (.Y(N3835), .A0(N3712), .A1(N4089), .B0(N4135), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I989 (.Y(N4033), .A0(N3712), .A1(N3382), .B0(N3450), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I990 (.Y(N3308), .A(N3712), .B(N2381));
AOI22XL cynw_cm_float_rcp_I991 (.Y(N3387), .A0(N3712), .A1(N3598), .B0(N3793), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I992 (.Y(N3593), .A0(N3712), .A1(N3584), .B0(N4132), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I993 (.Y(N3799), .A0(N3712), .A1(N3800), .B0(N3759), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I994 (.Y(N3996), .A0(N3712), .A1(N3392), .B0(N3838), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I995 (.Y(N3266), .A0(N3712), .A1(N3792), .B0(N3622), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I996 (.Y(N3475), .A0(N3712), .A1(N3792), .B0(N3520), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I997 (.Y(N3683), .A0(N3712), .A1(N3672), .B0(N3616), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I998 (.Y(N3882), .A0(N3712), .A1(N4074), .B0(N3382), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I999 (.Y(N4088), .A0(N3712), .A1(N3753), .B0(N3344), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1000 (.Y(N3358), .A0(N3712), .A1(N3838), .B0(N3393), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1001 (.Y(N3559), .A0(N3712), .A1(N3393), .B0(N3858), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1002 (.Y(N3766), .A0(N3712), .A1(N3974), .B0(N3828), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1003 (.Y(N3401), .A0(N3712), .A1(N3757), .B0(N3911), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1004 (.Y(N3611), .A0(N3712), .A1(N3938), .B0(N3467), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1005 (.Y(N3814), .A0(N3712), .A1(N3956), .B0(N3931), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1006 (.Y(N4012), .A0(N3712), .A1(N2381), .B0(N3616), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1007 (.Y(N3283), .A0(N3712), .A1(N3769), .B0(N3422), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1008 (.Y(N3491), .A0(N3712), .A1(a_man[18]), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1009 (.Y(N3695), .A0(N3712), .A1(N3446), .B0(N4030), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1010 (.Y(N3896), .A0(N3712), .A1(N3446), .B0(N3958), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1011 (.Y(N4104), .A0(N3712), .A1(N3974), .B0(N3240), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1012 (.Y(N3372), .A0(N3712), .A1(N4054), .B0(N3541), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1013 (.Y(N3572), .A0(N3712), .A1(N3639), .B0(N3967), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1014 (.Y(N3776), .A0(N3712), .A1(N3637), .B0(N3397), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1015 (.Y(N3977), .A0(N3712), .A1(N3492), .B0(N3524), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1016 (.Y(N3247), .A0(N3712), .A1(N3313), .B0(N3993), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1017 (.Y(N3453), .A0(N3712), .A1(N3889), .B0(N3258), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1018 (.Y(N3663), .A0(N3712), .A1(N3248), .B0(N3828), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1019 (.Y(N3862), .A(N3724), .B(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1020 (.Y(N3946), .A0(N3712), .A1(N3344), .B0(N3258), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1021 (.Y(N3214), .A0(N3712), .A1(a_man[17]), .B0(N3207), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1022 (.Y(N3416), .A0(N3712), .A1(N3533), .B0(N4089), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1023 (.Y(N3627), .A0(N3712), .A1(N2381), .B0(N3382), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I1024 (.Y(N3827), .A(N3712), .B(N2381));
NAND2XL cynw_cm_float_rcp_I1025 (.Y(N3330), .A(a_man[16]), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1026 (.Y(N3939), .A0(N3639), .A1(N3515), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1027 (.Y(N3905), .A0(N3639), .A1(N3721), .B0(N3342), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1028 (.Y(N3221), .A(N3639), .B(N3342));
AOI22XL cynw_cm_float_rcp_I1029 (.Y(N3836), .A0(N3639), .A1(N3220), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1030 (.Y(N3270), .A0(N3639), .A1(N3342), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1031 (.Y(N3360), .A0(N3639), .A1(N3342), .B0(N3220), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1032 (.Y(N3562), .A(N3639), .B(N3634));
AOI22XL cynw_cm_float_rcp_I1033 (.Y(N3235), .A0(N3639), .A1(N3867), .B0(N3480), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I1034 (.Y(N3442), .A(N3634), .B(a_man[18]));
NAND2XL cynw_cm_float_rcp_I1035 (.Y(N3603), .A(N3639), .B(N3634));
AOI22XL cynw_cm_float_rcp_I1036 (.Y(N4004), .A0(N3639), .A1(a_man[16]), .B0(N3721), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1037 (.Y(N3275), .A0(N3639), .A1(N3515), .B0(N3706), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1038 (.Y(N3483), .A(N3639), .B(N3480));
AOI22XL cynw_cm_float_rcp_I1039 (.Y(N4096), .A0(N3639), .A1(N3867), .B0(N3342), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1040 (.Y(N3789), .A0(N3639), .A1(N3721), .B0(N3515), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1041 (.Y(N4073), .A0(N3639), .A1(N3634), .B0(N3220), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1042 (.Y(N3223), .A0(N3639), .A1(N3342), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1043 (.Y(N3601), .A0(N3639), .A1(N3480), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1044 (.Y(N3273), .A0(N3639), .A1(N3867), .B0(N3750), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1045 (.Y(N3237), .A0(N3712), .A1(N3855), .B0(N3891), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1046 (.Y(N3444), .A0(N3712), .A1(N4024), .B0(N3548), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1047 (.Y(N3652), .A0(N3712), .A1(N3388), .B0(N4118), .B1(a_man[19]));
INVXL cynw_cm_float_rcp_I1048 (.Y(N3327), .A(N3486));
INVXL cynw_cm_float_rcp_I1049 (.Y(N3534), .A(N3299));
AOI22XL cynw_cm_float_rcp_I1050 (.Y(N3736), .A0(N3712), .A1(N3664), .B0(N3248), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1051 (.Y(N3701), .A0(N3712), .A1(N3603), .B0(N3330), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1052 (.Y(N3903), .A0(N3712), .A1(N4004), .B0(N3227), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1053 (.Y(N4110), .A0(N3712), .A1(N3275), .B0(N3939), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1054 (.Y(N3377), .A0(N3712), .A1(N3483), .B0(N3674), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1055 (.Y(N3576), .A0(N3712), .A1(N4096), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1056 (.Y(N3780), .A0(N3712), .A1(N3210), .B0(N3548), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1057 (.Y(N3981), .A0(N3712), .A1(N3956), .B0(N3464), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1058 (.Y(N3252), .A0(N3712), .A1(N3520), .B0(N3905), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1059 (.Y(N3457), .A0(N3712), .A1(N3221), .B0(N3874), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1060 (.Y(N3667), .A0(N3712), .A1(N4135), .B0(N3350), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1061 (.Y(N3866), .A0(N3712), .A1(N3450), .B0(N4099), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1062 (.Y(N4068), .A0(N3712), .A1(a_man[16]), .B0(N3806), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1063 (.Y(N3340), .A0(N3712), .A1(N3721), .B0(N3636), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1064 (.Y(N3748), .A0(N3712), .A1(N2381), .B0(N3641), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1065 (.Y(N3305), .A0(N3712), .A1(N3367), .B0(N3221), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1066 (.Y(N3512), .A0(N3712), .A1(N3789), .B0(N3836), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1067 (.Y(N3715), .A0(N3712), .A1(N3448), .B0(N3221), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1068 (.Y(N3919), .A0(N3712), .A1(N3623), .B0(N3315), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1069 (.Y(N4121), .A0(N3712), .A1(N4135), .B0(N3258), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1070 (.Y(N3385), .A0(N3712), .A1(N4073), .B0(N3277), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1071 (.Y(N3591), .A0(N3712), .A1(N3442), .B0(N3658), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1072 (.Y(N3797), .A0(N3712), .A1(N4115), .B0(N3854), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1073 (.Y(N3994), .A0(N3712), .A1(N3598), .B0(N3270), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1074 (.Y(N3264), .A0(N3712), .A1(N3223), .B0(N3240), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1075 (.Y(N3473), .A0(N3712), .A1(N3911), .B0(N3724), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1076 (.Y(N3681), .A0(N3712), .A1(N4089), .B0(N3360), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1077 (.Y(N3880), .A0(N3712), .A1(N3486), .B0(N3562), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1078 (.Y(N4086), .A0(N3712), .A1(N3791), .B0(N3235), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1079 (.Y(N3357), .A0(N3712), .A1(N3548), .B0(N3442), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1080 (.Y(N3557), .A0(N3712), .A1(N3442), .B0(N3258), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1081 (.Y(N3765), .A0(N3712), .A1(N3956), .B0(N3793), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1082 (.Y(N3966), .A0(N3712), .A1(N3601), .B0(a_man[18]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1083 (.Y(N3233), .A0(N3712), .A1(N3858), .B0(N3349), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1084 (.Y(N3438), .A0(N3712), .A1(N3524), .B0(N3874), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1085 (.Y(N3647), .A0(N3712), .A1(N3273), .B0(N3724), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1086 (.Y(N3847), .A0(N3712), .A1(N3639), .B0(N3641), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1087 (.Y(N3813), .A0(N3409), .A1(N3237), .B0(N3749), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1088 (.Y(N4011), .A0(N3409), .A1(N3444), .B0(N3951), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1089 (.Y(N3282), .A0(N3409), .A1(N3652), .B0(N3219), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1090 (.Y(N3490), .A0(N3409), .A1(N3344), .B0(N3424), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1091 (.Y(N3694), .A0(N3409), .A1(N3327), .B0(N3633), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1092 (.Y(N3895), .A0(N3409), .A1(N3534), .B0(N3835), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1093 (.Y(N4103), .A0(N3409), .A1(N3736), .B0(N4033), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1094 (.Y(N3371), .A0(N3409), .A1(N3709), .B0(N3308), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I1095 (.Y(N3571), .A(N3409), .B(N3709));
AOI22XL cynw_cm_float_rcp_I1096 (.Y(N3662), .A0(N3409), .A1(N3701), .B0(N3387), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1097 (.Y(N3861), .A0(N3409), .A1(N3903), .B0(N3593), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1098 (.Y(N4062), .A0(N3409), .A1(N4110), .B0(N3799), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1099 (.Y(N3336), .A0(N3409), .A1(N3377), .B0(N3996), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1100 (.Y(N3540), .A0(N3409), .A1(N3576), .B0(N3266), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1101 (.Y(N3744), .A0(N3409), .A1(N3780), .B0(N3475), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1102 (.Y(N3945), .A0(N3409), .A1(N3981), .B0(N3683), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1103 (.Y(N3213), .A0(N3409), .A1(N3252), .B0(N3882), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1104 (.Y(N3415), .A0(N3409), .A1(N3457), .B0(N4088), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1105 (.Y(N3626), .A0(N3409), .A1(N3667), .B0(N3358), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1106 (.Y(N3826), .A0(N3409), .A1(N3866), .B0(N3559), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1107 (.Y(N4025), .A0(N3409), .A1(N4068), .B0(N3766), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1108 (.Y(N3298), .A0(N3409), .A1(N3340), .B0(N3671), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1109 (.Y(N3506), .A0(N3409), .A1(N3445), .B0(N3870), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1110 (.Y(N3708), .A0(N3409), .A1(N3748), .B0(N3741), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1111 (.Y(N3913), .A0(N3409), .A1(N3926), .B0(N3741), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I1112 (.Y(N4117), .A(N3741), .B(a_man[20]));
NOR2XL cynw_cm_float_rcp_I1113 (.Y(N3587), .A(N3409), .B(N3558));
AOI22XL cynw_cm_float_rcp_I1114 (.Y(N3260), .A0(N3409), .A1(N3305), .B0(N3401), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1115 (.Y(N3466), .A0(N3409), .A1(N3512), .B0(N3611), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1116 (.Y(N3675), .A0(N3409), .A1(N3715), .B0(N3814), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1117 (.Y(N3873), .A0(N3409), .A1(N3919), .B0(N4012), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1118 (.Y(N4080), .A0(N3409), .A1(N4121), .B0(N3283), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1119 (.Y(N3348), .A0(N3409), .A1(N3385), .B0(N3491), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1120 (.Y(N3551), .A0(N3409), .A1(N3591), .B0(N3695), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1121 (.Y(N3758), .A0(N3409), .A1(N3797), .B0(N3896), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1122 (.Y(N3959), .A0(N3409), .A1(N3994), .B0(N4104), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1123 (.Y(N3226), .A0(N3409), .A1(N3264), .B0(N3372), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1124 (.Y(N3432), .A0(N3409), .A1(N3473), .B0(N3572), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1125 (.Y(N3640), .A0(N3409), .A1(N3681), .B0(N3776), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1126 (.Y(N3840), .A0(N3409), .A1(N3880), .B0(N3977), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1127 (.Y(N4043), .A0(N3409), .A1(N4086), .B0(N3247), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1128 (.Y(N3318), .A0(N3409), .A1(N3357), .B0(N3453), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1129 (.Y(N3523), .A0(N3409), .A1(N3557), .B0(N3663), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1130 (.Y(N3727), .A0(N3409), .A1(N3765), .B0(N3862), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1131 (.Y(N3930), .A0(N3409), .A1(N3966), .B0(N3536), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1132 (.Y(N4131), .A0(N3409), .A1(N3233), .B0(N3946), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1133 (.Y(N3396), .A0(N3409), .A1(N3438), .B0(N3214), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1134 (.Y(N3605), .A0(N3409), .A1(N3647), .B0(N3416), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1135 (.Y(N3807), .A0(N3409), .A1(N3847), .B0(N3627), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1136 (.Y(N4005), .A0(N3409), .A1(N3502), .B0(N3827), .B1(a_man[20]));
INVXL cynw_cm_float_rcp_I1137 (.Y(N4124), .A(N3750));
AOI22XL cynw_cm_float_rcp_I1138 (.Y(N3594), .A0(N3639), .A1(N3750), .B0(N3515), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1139 (.Y(N3997), .A0(N3639), .A1(a_man[17]), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1140 (.Y(N3731), .A0(N3639), .A1(a_man[17]), .B0(N3344), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1141 (.Y(N3402), .A0(N3639), .A1(a_man[16]), .B0(N3220), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1142 (.Y(N4106), .A0(N3639), .A1(N3342), .B0(N3706), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1143 (.Y(N4065), .A0(N3639), .A1(N3344), .B0(N3515), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1144 (.Y(N3291), .A0(N3639), .A1(N3515), .B0(N4034), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1145 (.Y(N4072), .A0(N3639), .A1(N4034), .B0(N3220), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1146 (.Y(N3599), .A0(N3639), .A1(N3634), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1147 (.Y(N3804), .A0(N3639), .A1(N3220), .B0(N3515), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1148 (.Y(N3287), .A0(N3712), .A1(N3990), .B0(N3317), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1149 (.Y(N3496), .A0(N3712), .A1(N3783), .B0(N4040), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1150 (.Y(N3699), .A0(N3712), .A1(N4044), .B0(N3429), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1151 (.Y(N3901), .A0(N3712), .A1(N3430), .B0(N3492), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1152 (.Y(N4109), .A0(N3712), .A1(N3417), .B0(N3990), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1153 (.Y(N3376), .A0(N3712), .A1(N4077), .B0(N3724), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1154 (.Y(N3575), .A0(N3712), .A1(N3691), .B0(N3388), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1155 (.Y(N3865), .A0(N3712), .A1(N4132), .B0(N4124), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1156 (.Y(N4066), .A0(N3712), .A1(N3492), .B0(N3588), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1157 (.Y(N3338), .A0(N3712), .A1(N3606), .B0(N3594), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1158 (.Y(N3543), .A0(N3712), .A1(N3291), .B0(N3608), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1159 (.Y(N3746), .A0(N3712), .A1(N4023), .B0(N3997), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1160 (.Y(N3949), .A0(N3712), .A1(N3606), .B0(N4042), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1161 (.Y(N3217), .A0(N3712), .A1(N3397), .B0(N3223), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1162 (.Y(N3421), .A0(N3712), .A1(N3395), .B0(N3546), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1163 (.Y(N3631), .A0(N3712), .A1(N3503), .B0(N3828), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1164 (.Y(N3832), .A0(N3712), .A1(N3297), .B0(N3825), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1165 (.Y(N4029), .A0(N3712), .A1(N3568), .B0(N3612), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1166 (.Y(N3303), .A0(N3712), .A1(N3492), .B0(N3315), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1167 (.Y(N3510), .A0(N3712), .A1(N3397), .B0(N3757), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1168 (.Y(N3713), .A0(N3712), .A1(N4072), .B0(N3612), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1169 (.Y(N3917), .A0(N3712), .A1(N3639), .B0(N3382), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1170 (.Y(N3471), .A0(N3712), .A1(N3297), .B0(N3731), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1171 (.Y(N3679), .A0(N3712), .A1(N3911), .B0(N3897), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1172 (.Y(N3878), .A0(N3712), .A1(N3246), .B0(N3911), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1173 (.Y(N4084), .A0(N3712), .A1(N3397), .B0(N3402), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1174 (.Y(N3354), .A0(N3712), .A1(N3429), .B0(N3722), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1175 (.Y(N3555), .A0(N3712), .A1(N4072), .B0(N3417), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1176 (.Y(N3763), .A0(N3712), .A1(N3858), .B0(N3623), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1177 (.Y(N3964), .A0(N3712), .A1(N3599), .B0(N4077), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1178 (.Y(N3231), .A0(N3712), .A1(N3804), .B0(N3267), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1179 (.Y(N3436), .A0(N3712), .A1(N3599), .B0(N4106), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1180 (.Y(N3645), .A0(N3712), .A1(N3838), .B0(N3809), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1181 (.Y(N3844), .A0(N3712), .A1(N3446), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1182 (.Y(N4048), .A0(N3712), .A1(N3225), .B0(N3897), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1183 (.Y(N3322), .A0(N3712), .A1(N4100), .B0(N3855), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1184 (.Y(N3529), .A0(N3712), .A1(N4106), .B0(N3672), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1185 (.Y(N3729), .A0(N3712), .A1(N4042), .B0(N4065), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1186 (.Y(N3933), .A0(N3712), .A1(N3769), .B0(N3927), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1187 (.Y(N4133), .A0(N3712), .A1(N3344), .B0(N3492), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1188 (.Y(N3398), .A0(N3712), .A1(N3486), .B0(N3524), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1189 (.Y(N3609), .A0(N3712), .A1(N3210), .B0(N3492), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1190 (.Y(N4009), .A0(N3712), .A1(N3382), .B0(N4118), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1191 (.Y(N3280), .A0(N3712), .A1(N3382), .B0(N4013), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1192 (.Y(N3274), .A(N3220), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1193 (.Y(N4053), .A0(N3639), .A1(N3515), .B0(N3721), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1194 (.Y(N3578), .A0(N3639), .A1(N3706), .B0(N3867), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1195 (.Y(N3782), .A0(N3639), .A1(N3342), .B0(N3344), .B1(a_man[18]));
NOR2XL cynw_cm_float_rcp_I1196 (.Y(N3341), .A(a_man[18]), .B(N3706));
AOI22XL cynw_cm_float_rcp_I1197 (.Y(N3307), .A0(N3639), .A1(N3867), .B0(N3463), .B1(a_man[18]));
NAND2XL cynw_cm_float_rcp_I1198 (.Y(N3514), .A(N3639), .B(N3480));
AOI22XL cynw_cm_float_rcp_I1199 (.Y(N4123), .A0(N3639), .A1(N3344), .B0(N3721), .B1(a_man[18]));
INVXL cynw_cm_float_rcp_I1200 (.Y(N3411), .A(N4034));
NAND2XL cynw_cm_float_rcp_I1201 (.Y(N3909), .A(N3480), .B(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1202 (.Y(N3655), .A0(N3639), .A1(N3220), .B0(N3634), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1203 (.Y(N3329), .A0(N3639), .A1(N3220), .B0(N3480), .B1(a_man[18]));
AOI22XL cynw_cm_float_rcp_I1204 (.Y(N3255), .A0(N3712), .A1(N3722), .B0(N3560), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1205 (.Y(N3459), .A0(N3712), .A1(N4100), .B0(N4065), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1206 (.Y(N3669), .A0(N3712), .A1(N3931), .B0(N3823), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1207 (.Y(N3869), .A0(N3712), .A1(N3524), .B0(N3388), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1208 (.Y(N4070), .A0(N3712), .A1(N3990), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1209 (.Y(N3343), .A0(N3712), .A1(N3492), .B0(N3486), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1210 (.Y(N3545), .A0(N3712), .A1(N3227), .B0(N3777), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1211 (.Y(N3751), .A0(N3712), .A1(N4013), .B0(N4135), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1212 (.Y(N4036), .A0(N3712), .A1(N3411), .B0(N3983), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1213 (.Y(N3310), .A0(N3712), .A1(N3990), .B0(N3274), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1214 (.Y(N3517), .A0(N3712), .A1(N4097), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1215 (.Y(N3718), .A0(N3712), .A1(N3578), .B0(N3330), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1216 (.Y(N3923), .A0(N3712), .A1(N3594), .B0(N3967), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1217 (.Y(N4126), .A(N3712), .B(N3993));
AOI22XL cynw_cm_float_rcp_I1218 (.Y(N3596), .A0(N3712), .A1(N3528), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1219 (.Y(N3802), .A0(N3712), .A1(N3909), .B0(N3752), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1220 (.Y(N3999), .A0(N3712), .A1(N3687), .B0(N4053), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1221 (.Y(N3269), .A0(N3712), .A1(N3931), .B0(N3921), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1222 (.Y(N3477), .A0(N3712), .A1(N3753), .B0(N3623), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1223 (.Y(N3685), .A0(N3712), .A1(N4071), .B0(N3721), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1224 (.Y(N3884), .A0(N3712), .A1(N3838), .B0(N3467), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1225 (.Y(N4091), .A0(N3712), .A1(a_man[17]), .B0(N4023), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1226 (.Y(N3359), .A0(N3712), .A1(a_man[18]), .B0(N3691), .B1(a_man[19]));
NAND2XL cynw_cm_float_rcp_I1227 (.Y(N3561), .A(N3664), .B(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1228 (.Y(N3441), .A0(N3712), .A1(N3674), .B0(N3731), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1229 (.Y(N3650), .A0(N3712), .A1(N3562), .B0(N4063), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1230 (.Y(N3851), .A0(N3712), .A1(N3563), .B0(N3578), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1231 (.Y(N4051), .A0(N3712), .A1(N3422), .B0(N3782), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1232 (.Y(N3326), .A0(N3712), .A1(N4078), .B0(N3349), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1233 (.Y(N3532), .A0(N3712), .A1(N3307), .B0(N4106), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1234 (.Y(N3733), .A0(N3712), .A1(N4044), .B0(N3350), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1235 (.Y(N3936), .A0(N3712), .A1(N3599), .B0(N3641), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1236 (.Y(N3204), .A0(N3712), .A1(N4054), .B0(N3608), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1237 (.Y(N3404), .A0(N3712), .A1(N3672), .B0(N3341), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1238 (.Y(N3615), .A0(N3712), .A1(N3854), .B0(N3872), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1239 (.Y(N3817), .A0(N3712), .A1(N4056), .B0(N3897), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1240 (.Y(N4016), .A0(N3712), .A1(N3655), .B0(N3440), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1241 (.Y(N3286), .A0(N3712), .A1(N3299), .B0(N3307), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1242 (.Y(N3495), .A0(N3712), .A1(N3350), .B0(N3514), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1243 (.Y(N3698), .A0(N3712), .A1(N3329), .B0(N3836), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1244 (.Y(N3900), .A0(N3712), .A1(N3562), .B0(N4123), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1245 (.Y(N4108), .A0(N3712), .A1(N4118), .B0(N3785), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I1246 (.Y(N3375), .A(N3712), .B(N3333));
AOI22XL cynw_cm_float_rcp_I1247 (.Y(N3980), .A0(N3712), .A1(N3344), .B0(N3838), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1248 (.Y(N3251), .A0(N3712), .A1(N3721), .B0(N3601), .B1(a_man[19]));
AOI22XL cynw_cm_float_rcp_I1249 (.Y(N3456), .A0(N3712), .A1(N3639), .B0(N3299), .B1(a_man[19]));
NOR2XL cynw_cm_float_rcp_I1250 (.Y(N3666), .A(N3712), .B(N3248));
AOI22XL cynw_cm_float_rcp_I1251 (.Y(N3420), .A0(N3409), .A1(N3255), .B0(N3287), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1252 (.Y(N3630), .A0(N3409), .A1(N3459), .B0(N3496), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1253 (.Y(N3831), .A0(N3409), .A1(N3669), .B0(N3699), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1254 (.Y(N4028), .A0(N3409), .A1(N3869), .B0(N3901), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1255 (.Y(N3302), .A0(N3409), .A1(N4070), .B0(N4109), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1256 (.Y(N3509), .A0(N3409), .A1(N3343), .B0(N3376), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1257 (.Y(N3711), .A0(N3409), .A1(N3545), .B0(N3575), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1258 (.Y(N3916), .A0(N3409), .A1(N3751), .B0(N3653), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1259 (.Y(N3992), .A0(N3409), .A1(N4036), .B0(N3865), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1260 (.Y(N3263), .A0(N3409), .A1(N3310), .B0(N4066), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1261 (.Y(N3470), .A0(N3409), .A1(N3517), .B0(N3338), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1262 (.Y(N3678), .A0(N3409), .A1(N3718), .B0(N3543), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1263 (.Y(N3877), .A0(N3409), .A1(N3923), .B0(N3746), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1264 (.Y(N4083), .A0(N3409), .A1(N4126), .B0(N3949), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1265 (.Y(N3353), .A0(N3409), .A1(N3596), .B0(N3217), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1266 (.Y(N3554), .A0(N3409), .A1(N3802), .B0(N3421), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1267 (.Y(N3762), .A0(N3409), .A1(N3999), .B0(N3631), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1268 (.Y(N3963), .A0(N3409), .A1(N3269), .B0(N3832), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1269 (.Y(N3230), .A0(N3409), .A1(N3477), .B0(N4029), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1270 (.Y(N3435), .A0(N3409), .A1(N3685), .B0(N3303), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1271 (.Y(N3644), .A0(N3409), .A1(N3884), .B0(N3510), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1272 (.Y(N3843), .A0(N3409), .A1(N4091), .B0(N3713), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1273 (.Y(N4047), .A0(N3409), .A1(N3359), .B0(N3917), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1274 (.Y(N3321), .A0(N3409), .A1(N3561), .B0(N3735), .B1(a_man[20]));
NOR2XL cynw_cm_float_rcp_I1275 (.Y(N3527), .A(N3409), .B(N4052));
AOI22XL cynw_cm_float_rcp_I1276 (.Y(N3607), .A0(N3409), .A1(N3441), .B0(N3471), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1277 (.Y(N3811), .A0(N3409), .A1(N3650), .B0(N3679), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1278 (.Y(N4008), .A0(N3409), .A1(N3851), .B0(N3878), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1279 (.Y(N3279), .A0(N3409), .A1(N4051), .B0(N4084), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1280 (.Y(N3489), .A0(N3409), .A1(N3326), .B0(N3354), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1281 (.Y(N3693), .A0(N3409), .A1(N3532), .B0(N3555), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1282 (.Y(N3893), .A0(N3409), .A1(N3733), .B0(N3763), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1283 (.Y(N4102), .A0(N3409), .A1(N3936), .B0(N3964), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1284 (.Y(N3370), .A0(N3409), .A1(N3204), .B0(N3231), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1285 (.Y(N3570), .A0(N3409), .A1(N3404), .B0(N3436), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1286 (.Y(N3775), .A0(N3409), .A1(N3615), .B0(N3645), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1287 (.Y(N3976), .A0(N3409), .A1(N3817), .B0(N3844), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1288 (.Y(N3245), .A0(N3409), .A1(N4016), .B0(N4048), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1289 (.Y(N3452), .A0(N3409), .A1(N3286), .B0(N3322), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1290 (.Y(N3661), .A0(N3409), .A1(N3495), .B0(N3529), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1291 (.Y(N3860), .A0(N3409), .A1(N3698), .B0(N3729), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1292 (.Y(N4061), .A0(N3409), .A1(N3900), .B0(N3933), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1293 (.Y(N3335), .A0(N3409), .A1(N4108), .B0(N4133), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1294 (.Y(N3539), .A0(N3409), .A1(N3375), .B0(N3398), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1295 (.Y(N3743), .A0(N3409), .A1(N3980), .B0(N3609), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1296 (.Y(N3944), .A0(N3409), .A1(N3251), .B0(N3671), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1297 (.Y(N3212), .A0(N3409), .A1(N3456), .B0(N4009), .B1(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1298 (.Y(N3414), .A0(N3409), .A1(N3666), .B0(N3280), .B1(a_man[20]));
NAND2XL cynw_cm_float_rcp_I1299 (.Y(N3625), .A(N3308), .B(a_man[20]));
AOI22XL cynw_cm_float_rcp_I1300 (.Y(N3505), .A0(N4112), .A1(N3420), .B0(N3813), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1301 (.Y(N3707), .A0(N4112), .A1(N3630), .B0(N4011), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1302 (.Y(N3912), .A0(N4112), .A1(N3831), .B0(N3282), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1303 (.Y(N4116), .A0(N4112), .A1(N4028), .B0(N3490), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1304 (.Y(N3383), .A0(N4112), .A1(N3302), .B0(N3694), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1305 (.Y(N3586), .A0(N4112), .A1(N3509), .B0(N3895), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1306 (.Y(N3794), .A0(N4112), .A1(N3711), .B0(N4103), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1307 (.Y(N3989), .A0(N4112), .A1(N3916), .B0(N3371), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1308 (.Y(N3259), .A0(N4112), .A1(N3864), .B0(N3571), .B1(a_man[21]));
NOR2XL cynw_cm_float_rcp_I1309 (.Y(N3400), .A(a_man[20]), .B(N3324));
NOR2XL cynw_cm_float_rcp_I1310 (.Y(N3465), .A(N3400), .B(N4112));
AOI22XL cynw_cm_float_rcp_I1311 (.Y(N4079), .A0(N4112), .A1(N3992), .B0(N3662), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1312 (.Y(N3347), .A0(N4112), .A1(N3263), .B0(N3861), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1313 (.Y(N3550), .A0(N4112), .A1(N3470), .B0(N4062), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1314 (.Y(N3756), .A0(N4112), .A1(N3678), .B0(N3336), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1315 (.Y(N3957), .A0(N4112), .A1(N3877), .B0(N3540), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1316 (.Y(N3224), .A0(N4112), .A1(N4083), .B0(N3744), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1317 (.Y(N3431), .A0(N4112), .A1(N3353), .B0(N3945), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1318 (.Y(N3638), .A0(N4112), .A1(N3554), .B0(N3213), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1319 (.Y(N3839), .A0(N4112), .A1(N3762), .B0(N3415), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1320 (.Y(N4041), .A0(N4112), .A1(N3963), .B0(N3626), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1321 (.Y(N3316), .A0(N4112), .A1(N3230), .B0(N3826), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1322 (.Y(N3522), .A0(N4112), .A1(N3435), .B0(N4025), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1323 (.Y(N3725), .A0(N4112), .A1(N3644), .B0(N3298), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1324 (.Y(N3928), .A0(N4112), .A1(N3843), .B0(N3506), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1325 (.Y(N4130), .A0(N4112), .A1(N4047), .B0(N3708), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1326 (.Y(N3394), .A0(N4112), .A1(N3321), .B0(N3913), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1327 (.Y(N3604), .A0(N4112), .A1(N3527), .B0(N4117), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1328 (.Y(N3276), .A0(N4112), .A1(N3607), .B0(N3260), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1329 (.Y(N3485), .A0(N4112), .A1(N3811), .B0(N3466), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1330 (.Y(N3690), .A0(N4112), .A1(N4008), .B0(N3675), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1331 (.Y(N3890), .A0(N4112), .A1(N3279), .B0(N3873), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1332 (.Y(N4098), .A0(N4112), .A1(N3489), .B0(N4080), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1333 (.Y(N3368), .A0(N4112), .A1(N3693), .B0(N3348), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1334 (.Y(N3567), .A0(N4112), .A1(N3893), .B0(N3551), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1335 (.Y(N3773), .A0(N4112), .A1(N4102), .B0(N3758), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1336 (.Y(N3973), .A0(N4112), .A1(N3370), .B0(N3959), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1337 (.Y(N3243), .A0(N4112), .A1(N3570), .B0(N3226), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1338 (.Y(N3449), .A0(N4112), .A1(N3775), .B0(N3432), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1339 (.Y(N3659), .A0(N4112), .A1(N3976), .B0(N3640), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1340 (.Y(N3857), .A0(N4112), .A1(N3245), .B0(N3840), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1341 (.Y(N4059), .A0(N4112), .A1(N3452), .B0(N4043), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1342 (.Y(N3332), .A0(N4112), .A1(N3661), .B0(N3318), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1343 (.Y(N3537), .A0(N4112), .A1(N3860), .B0(N3523), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1344 (.Y(N3740), .A0(N4112), .A1(N4061), .B0(N3727), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1345 (.Y(N3942), .A0(N4112), .A1(N3335), .B0(N3930), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1346 (.Y(N3208), .A0(N4112), .A1(N3539), .B0(N4131), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1347 (.Y(N3408), .A0(N4112), .A1(N3743), .B0(N3396), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1348 (.Y(N3620), .A0(N4112), .A1(N3944), .B0(N3605), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1349 (.Y(N3821), .A0(N4112), .A1(N3212), .B0(N3807), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1350 (.Y(N4021), .A0(N4112), .A1(N3414), .B0(N4005), .B1(a_man[21]));
AOI22XL cynw_cm_float_rcp_I1351 (.Y(N3294), .A0(N4112), .A1(N3625), .B0(N4069), .B1(a_man[21]));
INVX1 cynw_cm_float_rcp_I1352 (.Y(N3425), .A(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1353 (.Y(N449), .A0(N3425), .A1(N3505), .B0(N3216), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1354 (.Y(N450), .A0(N3425), .A1(N3707), .B0(N3419), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1355 (.Y(N451), .A0(N3425), .A1(N3912), .B0(N3629), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1356 (.Y(N452), .A0(N3425), .A1(N4116), .B0(N3830), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1357 (.Y(N453), .A0(N3425), .A1(N3383), .B0(N4027), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1358 (.Y(N454), .A0(N3425), .A1(N3586), .B0(N3301), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1359 (.Y(N455), .A0(N3425), .A1(N3794), .B0(N3508), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1360 (.Y(N456), .A0(N3425), .A1(N3989), .B0(N3915), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1361 (.Y(N457), .A0(N3425), .A1(N3259), .B0(N3590), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1363 (.Y(inst_cellmath__51[0]), .A0(N3425), .A1(N4079), .B0(N3262), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1364 (.Y(inst_cellmath__51[1]), .A0(N3425), .A1(N3347), .B0(N3469), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1365 (.Y(inst_cellmath__51[2]), .A0(N3425), .A1(N3550), .B0(N3677), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1366 (.Y(inst_cellmath__51[3]), .A0(N3425), .A1(N3756), .B0(N3876), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1367 (.Y(inst_cellmath__51[4]), .A0(N3425), .A1(N3957), .B0(N4082), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1368 (.Y(inst_cellmath__51[5]), .A0(N3425), .A1(N3224), .B0(N3352), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1369 (.Y(inst_cellmath__51[6]), .A0(N3425), .A1(N3431), .B0(N3553), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1370 (.Y(inst_cellmath__51[7]), .A0(N3425), .A1(N3638), .B0(N3761), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1371 (.Y(inst_cellmath__51[8]), .A0(N3425), .A1(N3839), .B0(N3962), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1372 (.Y(inst_cellmath__51[9]), .A0(N3425), .A1(N4041), .B0(N3229), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1373 (.Y(inst_cellmath__51[10]), .A0(N3425), .A1(N3316), .B0(N3434), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1374 (.Y(inst_cellmath__51[11]), .A0(N3425), .A1(N3522), .B0(N3643), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1375 (.Y(inst_cellmath__51[12]), .A0(N3425), .A1(N3725), .B0(N3842), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1376 (.Y(inst_cellmath__51[13]), .A0(N3425), .A1(N3928), .B0(N4046), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1377 (.Y(inst_cellmath__51[14]), .A0(N3425), .A1(N4130), .B0(N3320), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1378 (.Y(inst_cellmath__51[15]), .A0(N3425), .A1(N3394), .B0(N3526), .B1(a_man[22]));
NOR2XL cynw_cm_float_rcp_I1379 (.Y(inst_cellmath__51[16]), .A(a_man[22]), .B(N3604));
OAI2BB1X1 cynw_cm_float_rcp_I1380 (.Y(inst_cellmath__51[17]), .A0N(N3587), .A1N(a_man[21]), .B0(N3425));
AOI22XL cynw_cm_float_rcp_I1381 (.Y(N477), .A0(N3425), .A1(N3276), .B0(N3810), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1382 (.Y(N478), .A0(N3425), .A1(N3485), .B0(N4007), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1383 (.Y(N479), .A0(N3425), .A1(N3690), .B0(N3278), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1384 (.Y(N480), .A0(N3425), .A1(N3890), .B0(N3488), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1385 (.Y(N481), .A0(N3425), .A1(N4098), .B0(N3692), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1386 (.Y(N482), .A0(N3425), .A1(N3368), .B0(N3892), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1387 (.Y(N483), .A0(N3425), .A1(N3567), .B0(N4101), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1388 (.Y(N484), .A0(N3425), .A1(N3773), .B0(N3369), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1389 (.Y(N485), .A0(N3425), .A1(N3973), .B0(N3569), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1390 (.Y(N486), .A0(N3425), .A1(N3243), .B0(N3774), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1391 (.Y(N487), .A0(N3425), .A1(N3449), .B0(N3975), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1392 (.Y(N488), .A0(N3425), .A1(N3659), .B0(N3244), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1393 (.Y(N489), .A0(N3425), .A1(N3857), .B0(N3451), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1394 (.Y(N490), .A0(N3425), .A1(N4059), .B0(N3660), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1395 (.Y(N491), .A0(N3425), .A1(N3332), .B0(N3859), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1396 (.Y(N492), .A0(N3425), .A1(N3537), .B0(N4060), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1397 (.Y(N493), .A0(N3425), .A1(N3740), .B0(N3334), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1398 (.Y(N494), .A0(N3425), .A1(N3942), .B0(N3538), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1399 (.Y(N495), .A0(N3425), .A1(N3208), .B0(N3742), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1400 (.Y(N496), .A0(N3425), .A1(N3408), .B0(N3943), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1401 (.Y(N497), .A0(N3425), .A1(N3620), .B0(N3211), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1402 (.Y(N498), .A0(N3425), .A1(N3821), .B0(N3413), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1403 (.Y(N499), .A0(N3425), .A1(N4021), .B0(N3624), .B1(a_man[22]));
AOI22XL cynw_cm_float_rcp_I1404 (.Y(N500), .A0(N3425), .A1(N3294), .B0(N3824), .B1(a_man[22]));
NOR2XL cynw_cm_float_rcp_I1405 (.Y(N3894), .A(N4112), .B(N3952));
XOR2XL inst_cellmath__62_0_I4909 (.Y(N5380), .A(N2870), .B(N2652));
XOR2XL inst_cellmath__62_0_I4910 (.Y(N5115), .A(N2748), .B(N2794));
XOR2XL inst_cellmath__62_0_I4911 (.Y(N5186), .A(N2765), .B(N2610));
XOR2XL inst_cellmath__62_0_I4912 (.Y(N5259), .A(N2603), .B(N2751));
XOR2XL inst_cellmath__62_0_I4913 (.Y(N5334), .A(N2580), .B(N2892));
XOR2XL inst_cellmath__62_0_I4914 (.Y(N5072), .A(N2690), .B(N2710));
XOR2XL inst_cellmath__62_0_I4915 (.Y(N5146), .A(N2627), .B(N2851));
XOR2XL inst_cellmath__62_0_I4916 (.Y(N5219), .A(N2703), .B(N2667));
XOR2XL inst_cellmath__62_0_I4917 (.Y(N5292), .A(N2601), .B(N2812));
XOR2XL inst_cellmath__62_0_I4918 (.Y(N5365), .A(N2634), .B(N2625));
XOR2XL inst_cellmath__62_0_I4919 (.Y(N5101), .A(N2810), .B(N2768));
XOR2XL inst_cellmath__62_0_I4920 (.Y(N5174), .A(N2802), .B(N2588));
INVXL inst_cellmath__62_0_I1419 (.Y(N5246), .A(N449));
NOR2XL inst_cellmath__62_0_I1420 (.Y(inst_cellmath__62__W0[4]), .A(N5246), .B(N5380));
NOR2XL inst_cellmath__62_0_I1421 (.Y(inst_cellmath__62__W1[5]), .A(N5246), .B(N5115));
NOR2XL inst_cellmath__62_0_I1422 (.Y(N5156), .A(N5246), .B(N5186));
NOR2XL inst_cellmath__62_0_I1423 (.Y(N5300), .A(N5246), .B(N5259));
NOR2XL inst_cellmath__62_0_I1424 (.Y(N5110), .A(N5246), .B(N5334));
NOR2XL inst_cellmath__62_0_I1425 (.Y(N5256), .A(N5246), .B(N5072));
NOR2XL inst_cellmath__62_0_I1426 (.Y(N5067), .A(N5246), .B(N5146));
NOR2XL inst_cellmath__62_0_I1427 (.Y(N5214), .A(N5246), .B(N5219));
NOR2XL inst_cellmath__62_0_I1428 (.Y(N5363), .A(N5246), .B(N5292));
NOR2XL inst_cellmath__62_0_I1429 (.Y(N5172), .A(N5246), .B(N5365));
NOR2XL inst_cellmath__62_0_I1430 (.Y(N5318), .A(N5246), .B(N5101));
NOR2XL inst_cellmath__62_0_I1431 (.Y(N5127), .A(N5246), .B(N5174));
INVXL inst_cellmath__62_0_I1432 (.Y(N5322), .A(N450));
NOR2XL inst_cellmath__62_0_I1433 (.Y(inst_cellmath__62__W0[5]), .A(N5322), .B(N5380));
NOR2XL inst_cellmath__62_0_I1434 (.Y(inst_cellmath__62__W0[6]), .A(N5322), .B(N5115));
NOR2XL inst_cellmath__62_0_I1435 (.Y(N5367), .A(N5322), .B(N5186));
NOR2XL inst_cellmath__62_0_I1436 (.Y(N5176), .A(N5322), .B(N5259));
NOR2XL inst_cellmath__62_0_I1437 (.Y(N5325), .A(N5322), .B(N5334));
NOR2XL inst_cellmath__62_0_I1438 (.Y(N5134), .A(N5322), .B(N5072));
NOR2XL inst_cellmath__62_0_I1439 (.Y(N5280), .A(N5322), .B(N5146));
NOR2XL inst_cellmath__62_0_I1440 (.Y(N5089), .A(N5322), .B(N5219));
NOR2XL inst_cellmath__62_0_I1441 (.Y(N5236), .A(N5322), .B(N5292));
NOR2XL inst_cellmath__62_0_I1442 (.Y(N5386), .A(N5322), .B(N5365));
NOR2XL inst_cellmath__62_0_I1443 (.Y(N5195), .A(N5322), .B(N5101));
NOR2XL inst_cellmath__62_0_I1444 (.Y(N5340), .A(N5322), .B(N5174));
INVXL inst_cellmath__62_0_I1445 (.Y(N5397), .A(N451));
NOR2XL inst_cellmath__62_0_I1446 (.Y(N5287), .A(N5397), .B(N5380));
NOR2XL inst_cellmath__62_0_I1447 (.Y(N5095), .A(N5397), .B(N5115));
NOR2XL inst_cellmath__62_0_I1448 (.Y(N5241), .A(N5397), .B(N5186));
NOR2XL inst_cellmath__62_0_I1449 (.Y(N5391), .A(N5397), .B(N5259));
NOR2XL inst_cellmath__62_0_I1450 (.Y(N5199), .A(N5397), .B(N5334));
NOR2XL inst_cellmath__62_0_I1451 (.Y(N5346), .A(N5397), .B(N5072));
NOR2XL inst_cellmath__62_0_I1452 (.Y(N5158), .A(N5397), .B(N5146));
NOR2XL inst_cellmath__62_0_I1453 (.Y(N5304), .A(N5397), .B(N5219));
NOR2XL inst_cellmath__62_0_I1454 (.Y(N5114), .A(N5397), .B(N5292));
NOR2XL inst_cellmath__62_0_I1455 (.Y(N5260), .A(N5397), .B(N5365));
NOR2XL inst_cellmath__62_0_I1456 (.Y(N5071), .A(N5397), .B(N5101));
NOR2XL inst_cellmath__62_0_I1457 (.Y(N5218), .A(N5397), .B(N5174));
INVXL inst_cellmath__62_0_I1458 (.Y(N5132), .A(N452));
NOR2XL inst_cellmath__62_0_I1459 (.Y(N5163), .A(N5132), .B(N5380));
NOR2XL inst_cellmath__62_0_I1460 (.Y(N5309), .A(N5132), .B(N5115));
NOR2XL inst_cellmath__62_0_I1461 (.Y(N5120), .A(N5132), .B(N5186));
NOR2XL inst_cellmath__62_0_I1462 (.Y(N5265), .A(N5132), .B(N5259));
NOR2XL inst_cellmath__62_0_I1463 (.Y(N5076), .A(N5132), .B(N5334));
NOR2XL inst_cellmath__62_0_I1464 (.Y(N5224), .A(N5132), .B(N5072));
NOR2XL inst_cellmath__62_0_I1465 (.Y(N5372), .A(N5132), .B(N5146));
NOR2XL inst_cellmath__62_0_I1466 (.Y(N5179), .A(N5132), .B(N5219));
NOR2XL inst_cellmath__62_0_I1467 (.Y(N5328), .A(N5132), .B(N5292));
NOR2XL inst_cellmath__62_0_I1468 (.Y(N5139), .A(N5132), .B(N5365));
NOR2XL inst_cellmath__62_0_I1469 (.Y(N5284), .A(N5132), .B(N5101));
NOR2XL inst_cellmath__62_0_I1470 (.Y(N5092), .A(N5132), .B(N5174));
INVXL inst_cellmath__62_0_I1471 (.Y(N5205), .A(N453));
NOR2XL inst_cellmath__62_0_I1472 (.Y(N5379), .A(N5205), .B(N5380));
NOR2XL inst_cellmath__62_0_I1473 (.Y(N5185), .A(N5205), .B(N5115));
NOR2XL inst_cellmath__62_0_I1474 (.Y(N5333), .A(N5205), .B(N5186));
NOR2XL inst_cellmath__62_0_I1475 (.Y(N5145), .A(N5205), .B(N5259));
NOR2XL inst_cellmath__62_0_I1476 (.Y(N5291), .A(N5205), .B(N5334));
NOR2XL inst_cellmath__62_0_I1477 (.Y(N5099), .A(N5205), .B(N5072));
NOR2XL inst_cellmath__62_0_I1478 (.Y(N5245), .A(N5205), .B(N5146));
NOR2XL inst_cellmath__62_0_I1479 (.Y(N5396), .A(N5205), .B(N5219));
NOR2XL inst_cellmath__62_0_I1480 (.Y(N5204), .A(N5205), .B(N5292));
NOR2XL inst_cellmath__62_0_I1481 (.Y(N5353), .A(N5205), .B(N5365));
NOR2XL inst_cellmath__62_0_I1482 (.Y(N5162), .A(N5205), .B(N5101));
NOR2XL inst_cellmath__62_0_I1483 (.Y(N5308), .A(N5205), .B(N5174));
INVXL inst_cellmath__62_0_I1484 (.Y(N5278), .A(N454));
NOR2XL inst_cellmath__62_0_I1485 (.Y(N5249), .A(N5278), .B(N5380));
NOR2XL inst_cellmath__62_0_I1486 (.Y(N5401), .A(N5278), .B(N5115));
NOR2XL inst_cellmath__62_0_I1487 (.Y(N5208), .A(N5278), .B(N5186));
NOR2XL inst_cellmath__62_0_I1488 (.Y(N5358), .A(N5278), .B(N5259));
NOR2XL inst_cellmath__62_0_I1489 (.Y(N5166), .A(N5278), .B(N5334));
NOR2XL inst_cellmath__62_0_I1490 (.Y(N5312), .A(N5278), .B(N5072));
NOR2XL inst_cellmath__62_0_I1491 (.Y(N5122), .A(N5278), .B(N5146));
NOR2XL inst_cellmath__62_0_I1492 (.Y(N5268), .A(N5278), .B(N5219));
NOR2XL inst_cellmath__62_0_I1493 (.Y(N5079), .A(N5278), .B(N5292));
NOR2XL inst_cellmath__62_0_I1494 (.Y(N5229), .A(N5278), .B(N5365));
NOR2XL inst_cellmath__62_0_I1495 (.Y(N5377), .A(N5278), .B(N5101));
NOR2XL inst_cellmath__62_0_I1496 (.Y(N5183), .A(N5278), .B(N5174));
INVXL inst_cellmath__62_0_I1497 (.Y(N5355), .A(N455));
NOR2XL inst_cellmath__62_0_I1498 (.Y(N5129), .A(N5355), .B(N5380));
NOR2XL inst_cellmath__62_0_I1499 (.Y(N5274), .A(N5355), .B(N5115));
NOR2XL inst_cellmath__62_0_I1500 (.Y(N5083), .A(N5355), .B(N5186));
NOR2XL inst_cellmath__62_0_I1501 (.Y(N5231), .A(N5355), .B(N5259));
NOR2XL inst_cellmath__62_0_I1502 (.Y(N5382), .A(N5355), .B(N5334));
NOR2XL inst_cellmath__62_0_I1503 (.Y(N5189), .A(N5355), .B(N5072));
NOR2XL inst_cellmath__62_0_I1504 (.Y(N5337), .A(N5355), .B(N5146));
NOR2XL inst_cellmath__62_0_I1505 (.Y(N5148), .A(N5355), .B(N5219));
NOR2XL inst_cellmath__62_0_I1506 (.Y(N5295), .A(N5355), .B(N5292));
NOR2XL inst_cellmath__62_0_I1507 (.Y(N5104), .A(N5355), .B(N5365));
NOR2XL inst_cellmath__62_0_I1508 (.Y(N5247), .A(N5355), .B(N5101));
NOR2XL inst_cellmath__62_0_I1509 (.Y(N5399), .A(N5355), .B(N5174));
INVXL inst_cellmath__62_0_I1510 (.Y(N5086), .A(N456));
NOR2XL inst_cellmath__62_0_I1511 (.Y(N5342), .A(N5086), .B(N5380));
NOR2XL inst_cellmath__62_0_I1512 (.Y(N5154), .A(N5086), .B(N5115));
NOR2XL inst_cellmath__62_0_I1513 (.Y(N5299), .A(N5086), .B(N5186));
NOR2XL inst_cellmath__62_0_I1514 (.Y(N5108), .A(N5086), .B(N5259));
NOR2XL inst_cellmath__62_0_I1515 (.Y(N5254), .A(N5086), .B(N5334));
NOR2XL inst_cellmath__62_0_I1516 (.Y(N5066), .A(N5086), .B(N5072));
NOR2XL inst_cellmath__62_0_I1517 (.Y(N5212), .A(N5086), .B(N5146));
NOR2XL inst_cellmath__62_0_I1518 (.Y(N5361), .A(N5086), .B(N5219));
NOR2XL inst_cellmath__62_0_I1519 (.Y(N5171), .A(N5086), .B(N5292));
NOR2XL inst_cellmath__62_0_I1520 (.Y(N5316), .A(N5086), .B(N5365));
NOR2XL inst_cellmath__62_0_I1521 (.Y(N5125), .A(N5086), .B(N5101));
NOR2XL inst_cellmath__62_0_I1522 (.Y(N5272), .A(N5086), .B(N5174));
INVXL inst_cellmath__62_0_I1523 (.Y(N5164), .A(N457));
NOR2XL inst_cellmath__62_0_I1524 (.Y(N5220), .A(N5164), .B(N5380));
NOR2XL inst_cellmath__62_0_I1525 (.Y(N5366), .A(N5164), .B(N5115));
NOR2XL inst_cellmath__62_0_I1526 (.Y(N5175), .A(N5164), .B(N5186));
NOR2XL inst_cellmath__62_0_I1527 (.Y(N5323), .A(N5164), .B(N5259));
NOR2XL inst_cellmath__62_0_I1528 (.Y(N5133), .A(N5164), .B(N5334));
NOR2XL inst_cellmath__62_0_I1529 (.Y(N5279), .A(N5164), .B(N5072));
NOR2XL inst_cellmath__62_0_I1530 (.Y(N5087), .A(N5164), .B(N5146));
NOR2XL inst_cellmath__62_0_I1531 (.Y(N5235), .A(N5164), .B(N5219));
NOR2XL inst_cellmath__62_0_I1532 (.Y(N5385), .A(N5164), .B(N5292));
NOR2XL inst_cellmath__62_0_I1533 (.Y(N5193), .A(N5164), .B(N5365));
NOR2XL inst_cellmath__62_0_I1534 (.Y(N5339), .A(N5164), .B(N5101));
NOR2XL inst_cellmath__62_0_I1535 (.Y(N5152), .A(N5164), .B(N5174));
OR2XL inst_cellmath__62_0_I4921 (.Y(N5234), .A(a_man[22]), .B(N3465));
NOR2XL inst_cellmath__62_0_I1537 (.Y(N5094), .A(N5234), .B(N5380));
NOR2XL inst_cellmath__62_0_I1538 (.Y(N5240), .A(N5234), .B(N5115));
NOR2XL inst_cellmath__62_0_I1539 (.Y(N5389), .A(N5234), .B(N5186));
NOR2XL inst_cellmath__62_0_I1540 (.Y(N5198), .A(N5234), .B(N5259));
NOR2XL inst_cellmath__62_0_I1541 (.Y(N5345), .A(N5234), .B(N5334));
NOR2XL inst_cellmath__62_0_I1542 (.Y(N5157), .A(N5234), .B(N5072));
NOR2XL inst_cellmath__62_0_I1543 (.Y(N5303), .A(N5234), .B(N5146));
NOR2XL inst_cellmath__62_0_I1544 (.Y(N5113), .A(N5234), .B(N5219));
NOR2XL inst_cellmath__62_0_I1545 (.Y(N5258), .A(N5234), .B(N5292));
NOR2XL inst_cellmath__62_0_I1546 (.Y(N5070), .A(N5234), .B(N5365));
NOR2XL inst_cellmath__62_0_I1547 (.Y(N5217), .A(N5234), .B(N5101));
NOR2XL inst_cellmath__62_0_I1548 (.Y(inst_cellmath__62__W0[24]), .A(N5234), .B(N5174));
ADDHX1 inst_cellmath__62_0_I1549 (.CO(N5321), .S(inst_cellmath__62__W1[6]), .A(N5287), .B(N5156));
ADDHX1 inst_cellmath__62_0_I1550 (.CO(N5131), .S(inst_cellmath__62__W0[7]), .A(N5163), .B(N5300));
ADDFX1 inst_cellmath__62_0_I1551 (.CO(N5277), .S(inst_cellmath__62__W1[7]), .A(N5367), .B(N5095), .CI(N5321));
ADDHX1 inst_cellmath__62_0_I1552 (.CO(N5085), .S(N5354), .A(N5379), .B(N5176));
ADDFX1 inst_cellmath__62_0_I1553 (.CO(N5233), .S(inst_cellmath__62__W0[8]), .A(N5110), .B(N5309), .CI(N5241));
ADDFX1 inst_cellmath__62_0_I1554 (.CO(inst_cellmath__62__W0[9]), .S(inst_cellmath__62__W1[8]), .A(N5354), .B(N5131), .CI(N5277));
ADDHX1 inst_cellmath__62_0_I1555 (.CO(N5192), .S(N5119), .A(N5249), .B(N5391));
ADDFX1 inst_cellmath__62_0_I1556 (.CO(N5338), .S(N5264), .A(N5256), .B(N5185), .CI(N5120));
ADDFX1 inst_cellmath__62_0_I1557 (.CO(N5151), .S(N5075), .A(N5085), .B(N5325), .CI(N5119));
ADDFX1 inst_cellmath__62_0_I1558 (.CO(inst_cellmath__62__W0[10]), .S(inst_cellmath__62__W1[9]), .A(N5264), .B(N5233), .CI(N5075));
ADDHX1 inst_cellmath__62_0_I1559 (.CO(N5106), .S(N5371), .A(N5129), .B(N5265));
ADDFX1 inst_cellmath__62_0_I1560 (.CO(N5250), .S(N5178), .A(N5134), .B(N5401), .CI(N5333));
ADDFX1 inst_cellmath__62_0_I1561 (.CO(N5062), .S(N5327), .A(N5067), .B(N5199), .CI(N5192));
ADDFX1 inst_cellmath__62_0_I1562 (.CO(N5209), .S(N5138), .A(N5338), .B(N5371), .CI(N5178));
ADDFX1 inst_cellmath__62_0_I1563 (.CO(inst_cellmath__62__W0[11]), .S(inst_cellmath__62__W1[10]), .A(N5327), .B(N5151), .CI(N5138));
ADDHX1 inst_cellmath__62_0_I1564 (.CO(N5167), .S(N5091), .A(N5342), .B(N5145));
ADDFX1 inst_cellmath__62_0_I1565 (.CO(N5313), .S(N5238), .A(N5346), .B(N5274), .CI(N5208));
ADDFX1 inst_cellmath__62_0_I1566 (.CO(N5123), .S(N5388), .A(N5280), .B(N5076), .CI(N5214));
ADDFX1 inst_cellmath__62_0_I1567 (.CO(N5269), .S(N5197), .A(N5091), .B(N5106), .CI(N5250));
ADDFX1 inst_cellmath__62_0_I1568 (.CO(N5080), .S(N5344), .A(N5238), .B(N5062), .CI(N5388));
ADDFX1 inst_cellmath__62_0_I1569 (.CO(inst_cellmath__62__W0[12]), .S(inst_cellmath__62__W1[11]), .A(N5209), .B(N5197), .CI(N5344));
ADDHX1 inst_cellmath__62_0_I1570 (.CO(N5378), .S(N5302), .A(N5220), .B(N5358));
ADDFX1 inst_cellmath__62_0_I1571 (.CO(N5184), .S(N5112), .A(N5224), .B(N5154), .CI(N5083));
ADDFX1 inst_cellmath__62_0_I1572 (.CO(N5332), .S(N5257), .A(N5158), .B(N5291), .CI(N5363));
ADDFX1 inst_cellmath__62_0_I1573 (.CO(N5144), .S(N5069), .A(N5167), .B(N5089), .CI(N5302));
ADDFX1 inst_cellmath__62_0_I1574 (.CO(N5290), .S(N5216), .A(N5123), .B(N5313), .CI(N5112));
ADDFX1 inst_cellmath__62_0_I1575 (.CO(N5098), .S(N5364), .A(N5257), .B(N5269), .CI(N5069));
ADDFX1 inst_cellmath__62_0_I1576 (.CO(inst_cellmath__62__W0[13]), .S(inst_cellmath__62__W1[12]), .A(N5216), .B(N5080), .CI(N5364));
ADDHX1 inst_cellmath__62_0_I1577 (.CO(N5395), .S(N5320), .A(N5094), .B(N5231));
ADDFX1 inst_cellmath__62_0_I1578 (.CO(N5203), .S(N5130), .A(N5099), .B(N5366), .CI(N5299));
ADDFX1 inst_cellmath__62_0_I1579 (.CO(N5352), .S(N5276), .A(N5372), .B(N5166), .CI(N5236));
ADDFX1 inst_cellmath__62_0_I1580 (.CO(N5161), .S(N5084), .A(N5304), .B(N5172), .CI(N5378));
ADDFX1 inst_cellmath__62_0_I1581 (.CO(N5307), .S(N5232), .A(N5184), .B(N5320), .CI(N5332));
ADDFX1 inst_cellmath__62_0_I1582 (.CO(N5118), .S(N5384), .A(N5144), .B(N5130), .CI(N5276));
ADDFX1 inst_cellmath__62_0_I1583 (.CO(N5263), .S(N5190), .A(N5290), .B(N5084), .CI(N5232));
ADDFX1 inst_cellmath__62_0_I1584 (.CO(inst_cellmath__62__W0[14]), .S(inst_cellmath__62__W1[13]), .A(N5384), .B(N5098), .CI(N5190));
ADDFX1 inst_cellmath__62_0_I1585 (.CO(N5223), .S(N5150), .A(N5312), .B(N5240), .CI(N5175));
ADDFX1 inst_cellmath__62_0_I1586 (.CO(N5370), .S(N5296), .A(N5108), .B(N5382), .CI(N5245));
ADDFX1 inst_cellmath__62_0_I1587 (.CO(N5177), .S(N5105), .A(N5386), .B(N5114), .CI(N5179));
ADDFX1 inst_cellmath__62_0_I1588 (.CO(N5326), .S(N5248), .A(N5318), .B(N5395), .CI(N5203));
ADDFX1 inst_cellmath__62_0_I1589 (.CO(N5137), .S(N5400), .A(N5161), .B(N5352), .CI(N5150));
ADDFX1 inst_cellmath__62_0_I1590 (.CO(N5283), .S(N5207), .A(N5105), .B(N5296), .CI(N5307));
ADDFX1 inst_cellmath__62_0_I1591 (.CO(N5090), .S(N5357), .A(N5118), .B(N5248), .CI(N5400));
ADDFX1 inst_cellmath__62_0_I1592 (.CO(inst_cellmath__62__W0[15]), .S(inst_cellmath__62__W1[14]), .A(N5263), .B(N5207), .CI(N5357));
ADDFX1 inst_cellmath__62_0_I1593 (.CO(N5387), .S(N5311), .A(N5254), .B(N5189), .CI(N5323));
ADDFX1 inst_cellmath__62_0_I1594 (.CO(N5196), .S(N5121), .A(N5122), .B(N5389), .CI(N5328));
ADDFX1 inst_cellmath__62_0_I1595 (.CO(N5343), .S(N5267), .A(N5396), .B(N5260), .CI(N5195));
ADDFX1 inst_cellmath__62_0_I1596 (.CO(N5155), .S(N5078), .A(N5223), .B(N5127), .CI(N5370));
ADDFX1 inst_cellmath__62_0_I1597 (.CO(N5301), .S(N5228), .A(N5311), .B(N5177), .CI(N5326));
ADDFX1 inst_cellmath__62_0_I1598 (.CO(N5111), .S(N5376), .A(N5267), .B(N5121), .CI(N5137));
ADDFX1 inst_cellmath__62_0_I1599 (.CO(N5255), .S(N5182), .A(N5283), .B(N5078), .CI(N5228));
ADDFX1 inst_cellmath__62_0_I1600 (.CO(inst_cellmath__62__W0[16]), .S(inst_cellmath__62__W1[15]), .A(N5376), .B(N5090), .CI(N5182));
ADDHX1 inst_cellmath__62_0_I1601 (.CO(N5215), .S(N5143), .A(N5066), .B(N5337));
ADDFX1 inst_cellmath__62_0_I1602 (.CO(N5362), .S(N5289), .A(N5198), .B(N5133), .CI(N5204));
ADDFX1 inst_cellmath__62_0_I1603 (.CO(N5173), .S(N5097), .A(N5268), .B(N5139), .CI(N5071));
ADDFX1 inst_cellmath__62_0_I1604 (.CO(N5319), .S(N5244), .A(N5143), .B(N5340), .CI(N5387));
ADDFX1 inst_cellmath__62_0_I1605 (.CO(N5126), .S(N5393), .A(N5343), .B(N5196), .CI(N5289));
ADDFX1 inst_cellmath__62_0_I1606 (.CO(N5273), .S(N5201), .A(N5097), .B(N5155), .CI(N5244));
ADDFX1 inst_cellmath__62_0_I1607 (.CO(N5081), .S(N5349), .A(N5393), .B(N5301), .CI(N5111));
ADDFX1 inst_cellmath__62_0_I1608 (.CO(inst_cellmath__62__W0[17]), .S(inst_cellmath__62__W1[16]), .A(N5255), .B(N5201), .CI(N5349));
ADDFX1 inst_cellmath__62_0_I1609 (.CO(N5381), .S(N5305), .A(N5345), .B(N5279), .CI(N5212));
ADDFX1 inst_cellmath__62_0_I1610 (.CO(N5187), .S(N5116), .A(N5353), .B(N5079), .CI(N5148));
ADDFX1 inst_cellmath__62_0_I1611 (.CO(N5335), .S(N5261), .A(N5218), .B(N5284), .CI(N5215));
ADDFX1 inst_cellmath__62_0_I1612 (.CO(N5147), .S(N5073), .A(N5173), .B(N5362), .CI(N5305));
ADDFX1 inst_cellmath__62_0_I1613 (.CO(N5293), .S(N5221), .A(N5116), .B(N5319), .CI(N5261));
ADDFX1 inst_cellmath__62_0_I1614 (.CO(N5102), .S(N5368), .A(N5073), .B(N5126), .CI(N5273));
ADDFX1 inst_cellmath__62_0_I1615 (.CO(inst_cellmath__62__W0[18]), .S(inst_cellmath__62__W1[17]), .A(N5081), .B(N5221), .CI(N5368));
ADDFX1 inst_cellmath__62_0_I1616 (.CO(N5398), .S(N5324), .A(N5087), .B(N5157), .CI(N5295));
ADDFX1 inst_cellmath__62_0_I1617 (.CO(N5206), .S(N5135), .A(N5361), .B(N5229), .CI(N5162));
ADDFX1 inst_cellmath__62_0_I1618 (.CO(N5356), .S(N5281), .A(N5381), .B(N5092), .CI(N5187));
ADDFX1 inst_cellmath__62_0_I1619 (.CO(N5165), .S(N5088), .A(N5324), .B(N5335), .CI(N5135));
ADDFX1 inst_cellmath__62_0_I1620 (.CO(N5310), .S(N5237), .A(N5281), .B(N5147), .CI(N5293));
ADDFX1 inst_cellmath__62_0_I1621 (.CO(inst_cellmath__62__W0[19]), .S(inst_cellmath__62__W1[18]), .A(N5102), .B(N5088), .CI(N5237));
ADDFX1 inst_cellmath__62_0_I1622 (.CO(N5266), .S(N5194), .A(N5171), .B(N5303), .CI(N5235));
ADDFX1 inst_cellmath__62_0_I1623 (.CO(N5077), .S(N5341), .A(N5377), .B(N5104), .CI(N5308));
ADDFX1 inst_cellmath__62_0_I1624 (.CO(N5226), .S(N5153), .A(N5206), .B(N5398), .CI(N5194));
ADDFX1 inst_cellmath__62_0_I1625 (.CO(N5374), .S(N5297), .A(N5356), .B(N5341), .CI(N5165));
ADDFX1 inst_cellmath__62_0_I1626 (.CO(inst_cellmath__62__W0[20]), .S(inst_cellmath__62__W1[19]), .A(N5310), .B(N5153), .CI(N5297));
ADDFX1 inst_cellmath__62_0_I1627 (.CO(N5330), .S(N5252), .A(N5316), .B(N5385), .CI(N5113));
ADDFX1 inst_cellmath__62_0_I1628 (.CO(N5141), .S(N5064), .A(N5183), .B(N5247), .CI(N5266));
ADDFX1 inst_cellmath__62_0_I1629 (.CO(N5286), .S(N5211), .A(N5252), .B(N5077), .CI(N5064));
ADDFX1 inst_cellmath__62_0_I1630 (.CO(inst_cellmath__62__W0[21]), .S(inst_cellmath__62__W1[20]), .A(N5374), .B(N5226), .CI(N5211));
ADDFX1 inst_cellmath__62_0_I1631 (.CO(N5242), .S(N5169), .A(N5193), .B(N5258), .CI(N5125));
ADDFX1 inst_cellmath__62_0_I1632 (.CO(N5390), .S(N5315), .A(N5330), .B(N5399), .CI(N5169));
ADDFX1 inst_cellmath__62_0_I1633 (.CO(inst_cellmath__62__W1[22]), .S(inst_cellmath__62__W1[21]), .A(N5315), .B(N5141), .CI(N5286));
ADDFX1 inst_cellmath__62_0_I1634 (.CO(N5347), .S(N5270), .A(N5339), .B(N5070), .CI(N5272));
ADDFX1 inst_cellmath__62_0_I1635 (.CO(inst_cellmath__62__W1[23]), .S(inst_cellmath__62__W0[22]), .A(N5270), .B(N5242), .CI(N5390));
ADDFX1 inst_cellmath__62_0_I1636 (.CO(inst_cellmath__62__W1[24]), .S(inst_cellmath__62__W0[23]), .A(N5152), .B(N5217), .CI(N5347));
INVXL inst_cellmath__63_0_I1637 (.Y(N6075), .A(inst_cellmath__51[0]));
INVXL inst_cellmath__63_0_I1638 (.Y(N6531), .A(inst_cellmath__51[1]));
INVXL inst_cellmath__63_0_I1639 (.Y(N6120), .A(inst_cellmath__51[2]));
INVXL inst_cellmath__63_0_I1640 (.Y(N6576), .A(inst_cellmath__51[3]));
INVXL inst_cellmath__63_0_I1641 (.Y(N6166), .A(inst_cellmath__51[4]));
INVXL inst_cellmath__63_0_I1642 (.Y(N5759), .A(inst_cellmath__51[5]));
INVXL inst_cellmath__63_0_I1643 (.Y(N6215), .A(inst_cellmath__51[6]));
INVXL inst_cellmath__63_0_I1644 (.Y(N5808), .A(inst_cellmath__51[7]));
INVXL inst_cellmath__63_0_I1645 (.Y(N6258), .A(inst_cellmath__51[8]));
INVXL inst_cellmath__63_0_I1646 (.Y(N5850), .A(inst_cellmath__51[9]));
INVXL inst_cellmath__63_0_I1647 (.Y(N6303), .A(inst_cellmath__51[10]));
INVXL inst_cellmath__63_0_I1648 (.Y(N5895), .A(inst_cellmath__51[11]));
INVXL inst_cellmath__63_0_I1649 (.Y(N6354), .A(inst_cellmath__51[12]));
INVXL inst_cellmath__63_0_I1650 (.Y(N5945), .A(inst_cellmath__51[13]));
INVXL inst_cellmath__63_0_I1651 (.Y(N6401), .A(inst_cellmath__51[14]));
INVXL inst_cellmath__63_0_I1652 (.Y(N5990), .A(inst_cellmath__51[15]));
INVXL inst_cellmath__63_0_I1653 (.Y(N6444), .A(inst_cellmath__51[16]));
INVXL inst_cellmath__63_0_I1654 (.Y(N6033), .A(inst_cellmath__51[17]));
INVXL inst_cellmath__63_0_I1655 (.Y(N6299), .A(a_man[0]));
NOR2XL inst_cellmath__63_0_I1658 (.Y(N5969), .A(N6299), .B(N6120));
NOR2XL inst_cellmath__63_0_I1659 (.Y(N6347), .A(N6299), .B(N6576));
NOR2XL inst_cellmath__63_0_I1660 (.Y(N5859), .A(N6299), .B(N6166));
NOR2XL inst_cellmath__63_0_I1661 (.Y(N6232), .A(N6299), .B(N5759));
NOR2XL inst_cellmath__63_0_I1662 (.Y(N5748), .A(N6299), .B(N6215));
NOR2XL inst_cellmath__63_0_I1663 (.Y(N6126), .A(N6299), .B(N5808));
NOR2XL inst_cellmath__63_0_I1664 (.Y(N6501), .A(N6299), .B(N6258));
NOR2XL inst_cellmath__63_0_I1665 (.Y(N6016), .A(N6299), .B(N5850));
NOR2XL inst_cellmath__63_0_I1666 (.Y(N6396), .A(N6299), .B(N6303));
NOR2XL inst_cellmath__63_0_I1667 (.Y(N5904), .A(N6299), .B(N5895));
NOR2XL inst_cellmath__63_0_I1668 (.Y(N6280), .A(N6299), .B(N6354));
NOR2XL inst_cellmath__63_0_I1669 (.Y(N5797), .A(N6299), .B(N5945));
NOR2XL inst_cellmath__63_0_I1670 (.Y(N6170), .A(N6299), .B(N6401));
NOR2XL inst_cellmath__63_0_I1671 (.Y(N6548), .A(N6299), .B(N5990));
NOR2XL inst_cellmath__63_0_I1672 (.Y(N6060), .A(N6299), .B(N6444));
NOR2XL inst_cellmath__63_0_I1673 (.Y(N6436), .A(N6299), .B(N6033));
INVXL inst_cellmath__63_0_I1674 (.Y(N6568), .A(a_man[1]));
NOR2XL inst_cellmath__63_0_I1676 (.Y(inst_cellmath__63__W0[2]), .A(N6568), .B(N6531));
NOR2XL inst_cellmath__63_0_I1677 (.Y(N6377), .A(N6568), .B(N6120));
NOR2XL inst_cellmath__63_0_I1678 (.Y(N5887), .A(N6568), .B(N6576));
NOR2XL inst_cellmath__63_0_I1679 (.Y(N6263), .A(N6568), .B(N6166));
NOR2XL inst_cellmath__63_0_I1680 (.Y(N5779), .A(N6568), .B(N5759));
NOR2XL inst_cellmath__63_0_I1681 (.Y(N6152), .A(N6568), .B(N6215));
NOR2XL inst_cellmath__63_0_I1682 (.Y(N6533), .A(N6568), .B(N5808));
NOR2XL inst_cellmath__63_0_I1683 (.Y(N6040), .A(N6568), .B(N6258));
NOR2XL inst_cellmath__63_0_I1684 (.Y(N6420), .A(N6568), .B(N5850));
NOR2XL inst_cellmath__63_0_I1685 (.Y(N5933), .A(N6568), .B(N6303));
NOR2XL inst_cellmath__63_0_I1686 (.Y(N6309), .A(N6568), .B(N5895));
NOR2XL inst_cellmath__63_0_I1687 (.Y(N5824), .A(N6568), .B(N6354));
NOR2XL inst_cellmath__63_0_I1688 (.Y(N6199), .A(N6568), .B(N5945));
NOR2XL inst_cellmath__63_0_I1689 (.Y(N6578), .A(N6568), .B(N6401));
NOR2XL inst_cellmath__63_0_I1690 (.Y(N6086), .A(N6568), .B(N5990));
NOR2XL inst_cellmath__63_0_I1691 (.Y(N6467), .A(N6568), .B(N6444));
NOR2XL inst_cellmath__63_0_I1692 (.Y(N5980), .A(N6568), .B(N6033));
INVXL inst_cellmath__63_0_I1693 (.Y(N5973), .A(a_man[2]));
NOR2XL inst_cellmath__63_0_I1694 (.Y(N6027), .A(N5973), .B(N6075));
NOR2XL inst_cellmath__63_0_I1695 (.Y(N6406), .A(N5973), .B(N6531));
NOR2XL inst_cellmath__63_0_I1696 (.Y(N5916), .A(N5973), .B(N6120));
NOR2XL inst_cellmath__63_0_I1697 (.Y(N6291), .A(N5973), .B(N6576));
NOR2XL inst_cellmath__63_0_I1698 (.Y(N5809), .A(N5973), .B(N6166));
NOR2XL inst_cellmath__63_0_I1699 (.Y(N6184), .A(N5973), .B(N5759));
NOR2XL inst_cellmath__63_0_I1700 (.Y(N6558), .A(N5973), .B(N6215));
NOR2XL inst_cellmath__63_0_I1701 (.Y(N6071), .A(N5973), .B(N5808));
NOR2XL inst_cellmath__63_0_I1702 (.Y(N6450), .A(N5973), .B(N6258));
NOR2XL inst_cellmath__63_0_I1703 (.Y(N5962), .A(N5973), .B(N5850));
NOR2XL inst_cellmath__63_0_I1704 (.Y(N6339), .A(N5973), .B(N6303));
NOR2XL inst_cellmath__63_0_I1705 (.Y(N5851), .A(N5973), .B(N5895));
NOR2XL inst_cellmath__63_0_I1706 (.Y(N6225), .A(N5973), .B(N6354));
NOR2XL inst_cellmath__63_0_I1707 (.Y(N5741), .A(N5973), .B(N5945));
NOR2XL inst_cellmath__63_0_I1708 (.Y(N6116), .A(N5973), .B(N6401));
NOR2XL inst_cellmath__63_0_I1709 (.Y(N6492), .A(N5973), .B(N5990));
NOR2XL inst_cellmath__63_0_I1710 (.Y(N6007), .A(N5973), .B(N6444));
NOR2XL inst_cellmath__63_0_I1711 (.Y(N6387), .A(N5973), .B(N6033));
NOR2XL inst_cellmath__63_0_I1713 (.Y(N6430), .A(N2875), .B(N6075));
NOR2XL inst_cellmath__63_0_I1714 (.Y(N5947), .A(N2875), .B(N6531));
NOR2XL inst_cellmath__63_0_I1715 (.Y(N6323), .A(N2875), .B(N6120));
NOR2XL inst_cellmath__63_0_I1716 (.Y(N5836), .A(N2875), .B(N6576));
NOR2XL inst_cellmath__63_0_I1717 (.Y(N6211), .A(N2875), .B(N6166));
NOR2XL inst_cellmath__63_0_I1718 (.Y(N5728), .A(N2875), .B(N5759));
NOR2XL inst_cellmath__63_0_I1719 (.Y(N6098), .A(N2875), .B(N6215));
NOR2XL inst_cellmath__63_0_I1720 (.Y(N6479), .A(N2875), .B(N5808));
NOR2XL inst_cellmath__63_0_I1721 (.Y(N5992), .A(N2875), .B(N6258));
NOR2XL inst_cellmath__63_0_I1722 (.Y(N6367), .A(N2875), .B(N5850));
NOR2XL inst_cellmath__63_0_I1723 (.Y(N5879), .A(N2875), .B(N6303));
NOR2XL inst_cellmath__63_0_I1724 (.Y(N6254), .A(N2875), .B(N5895));
NOR2XL inst_cellmath__63_0_I1725 (.Y(N5769), .A(N2875), .B(N6354));
NOR2XL inst_cellmath__63_0_I1726 (.Y(N6144), .A(N2875), .B(N5945));
NOR2XL inst_cellmath__63_0_I1727 (.Y(N6523), .A(N2875), .B(N6401));
NOR2XL inst_cellmath__63_0_I1728 (.Y(N6032), .A(N2875), .B(N5990));
NOR2XL inst_cellmath__63_0_I1729 (.Y(N6412), .A(N2875), .B(N6444));
NOR2XL inst_cellmath__63_0_I1730 (.Y(N5927), .A(N2875), .B(N6033));
NOR2XL inst_cellmath__63_0_I1732 (.Y(N5975), .A(N2631), .B(N6075));
NOR2XL inst_cellmath__63_0_I1733 (.Y(N6351), .A(N2631), .B(N6531));
NOR2XL inst_cellmath__63_0_I1734 (.Y(N5863), .A(N2631), .B(N6120));
NOR2XL inst_cellmath__63_0_I1735 (.Y(N6238), .A(N2631), .B(N6576));
NOR2XL inst_cellmath__63_0_I1736 (.Y(N5752), .A(N2631), .B(N6166));
NOR2XL inst_cellmath__63_0_I1737 (.Y(N6130), .A(N2631), .B(N5759));
NOR2XL inst_cellmath__63_0_I1738 (.Y(N6507), .A(N2631), .B(N6215));
NOR2XL inst_cellmath__63_0_I1739 (.Y(N6020), .A(N2631), .B(N5808));
NOR2XL inst_cellmath__63_0_I1740 (.Y(N6398), .A(N2631), .B(N6258));
NOR2XL inst_cellmath__63_0_I1741 (.Y(N5910), .A(N2631), .B(N5850));
NOR2XL inst_cellmath__63_0_I1742 (.Y(N6283), .A(N2631), .B(N6303));
NOR2XL inst_cellmath__63_0_I1743 (.Y(N5800), .A(N2631), .B(N5895));
NOR2XL inst_cellmath__63_0_I1744 (.Y(N6175), .A(N2631), .B(N6354));
NOR2XL inst_cellmath__63_0_I1745 (.Y(N6551), .A(N2631), .B(N5945));
NOR2XL inst_cellmath__63_0_I1746 (.Y(N6063), .A(N2631), .B(N6401));
NOR2XL inst_cellmath__63_0_I1747 (.Y(N6440), .A(N2631), .B(N5990));
NOR2XL inst_cellmath__63_0_I1748 (.Y(N5954), .A(N2631), .B(N6444));
NOR2XL inst_cellmath__63_0_I1749 (.Y(N6331), .A(N2631), .B(N6033));
NOR2XL inst_cellmath__63_0_I1751 (.Y(N6381), .A(N2698), .B(N6075));
NOR2XL inst_cellmath__63_0_I1752 (.Y(N5890), .A(N2698), .B(N6531));
NOR2XL inst_cellmath__63_0_I1753 (.Y(N6266), .A(N2698), .B(N6120));
NOR2XL inst_cellmath__63_0_I1754 (.Y(N5783), .A(N2698), .B(N6576));
NOR2XL inst_cellmath__63_0_I1755 (.Y(N6155), .A(N2698), .B(N6166));
NOR2XL inst_cellmath__63_0_I1756 (.Y(N6536), .A(N2698), .B(N5759));
NOR2XL inst_cellmath__63_0_I1757 (.Y(N6045), .A(N2698), .B(N6215));
NOR2XL inst_cellmath__63_0_I1758 (.Y(N6422), .A(N2698), .B(N5808));
NOR2XL inst_cellmath__63_0_I1759 (.Y(N5937), .A(N2698), .B(N6258));
NOR2XL inst_cellmath__63_0_I1760 (.Y(N6314), .A(N2698), .B(N5850));
NOR2XL inst_cellmath__63_0_I1761 (.Y(N5828), .A(N2698), .B(N6303));
NOR2XL inst_cellmath__63_0_I1762 (.Y(N6203), .A(N2698), .B(N5895));
NOR2XL inst_cellmath__63_0_I1763 (.Y(N5722), .A(N2698), .B(N6354));
NOR2XL inst_cellmath__63_0_I1764 (.Y(N6090), .A(N2698), .B(N5945));
NOR2XL inst_cellmath__63_0_I1765 (.Y(N6471), .A(N2698), .B(N6401));
NOR2XL inst_cellmath__63_0_I1766 (.Y(N5983), .A(N2698), .B(N5990));
NOR2XL inst_cellmath__63_0_I1767 (.Y(N6359), .A(N2698), .B(N6444));
NOR2XL inst_cellmath__63_0_I1768 (.Y(N5871), .A(N2698), .B(N6033));
NOR2XL inst_cellmath__63_0_I1770 (.Y(N5919), .A(N2772), .B(N6075));
NOR2XL inst_cellmath__63_0_I1771 (.Y(N6293), .A(N2772), .B(N6531));
NOR2XL inst_cellmath__63_0_I1772 (.Y(N5811), .A(N2772), .B(N6120));
NOR2XL inst_cellmath__63_0_I1773 (.Y(N6187), .A(N2772), .B(N6576));
NOR2XL inst_cellmath__63_0_I1774 (.Y(N6560), .A(N2772), .B(N6166));
NOR2XL inst_cellmath__63_0_I1775 (.Y(N6074), .A(N2772), .B(N5759));
NOR2XL inst_cellmath__63_0_I1776 (.Y(N6453), .A(N2772), .B(N6215));
NOR2XL inst_cellmath__63_0_I1777 (.Y(N5964), .A(N2772), .B(N5808));
NOR2XL inst_cellmath__63_0_I1778 (.Y(N6342), .A(N2772), .B(N6258));
NOR2XL inst_cellmath__63_0_I1779 (.Y(N5854), .A(N2772), .B(N5850));
NOR2XL inst_cellmath__63_0_I1780 (.Y(N6227), .A(N2772), .B(N6303));
NOR2XL inst_cellmath__63_0_I1781 (.Y(N5743), .A(N2772), .B(N5895));
NOR2XL inst_cellmath__63_0_I1782 (.Y(N6119), .A(N2772), .B(N6354));
NOR2XL inst_cellmath__63_0_I1783 (.Y(N6495), .A(N2772), .B(N5945));
NOR2XL inst_cellmath__63_0_I1784 (.Y(N6010), .A(N2772), .B(N6401));
NOR2XL inst_cellmath__63_0_I1785 (.Y(N6390), .A(N2772), .B(N5990));
NOR2XL inst_cellmath__63_0_I1786 (.Y(N5898), .A(N2772), .B(N6444));
NOR2XL inst_cellmath__63_0_I1787 (.Y(N6274), .A(N2772), .B(N6033));
NOR2XL inst_cellmath__63_0_I1789 (.Y(N6326), .A(N2579), .B(N6075));
NOR2XL inst_cellmath__63_0_I1790 (.Y(N5839), .A(N2579), .B(N6531));
NOR2XL inst_cellmath__63_0_I1791 (.Y(N6214), .A(N2579), .B(N6120));
NOR2XL inst_cellmath__63_0_I1792 (.Y(N5731), .A(N2579), .B(N6576));
NOR2XL inst_cellmath__63_0_I1793 (.Y(N6101), .A(N2579), .B(N6166));
NOR2XL inst_cellmath__63_0_I1794 (.Y(N6482), .A(N2579), .B(N5759));
NOR2XL inst_cellmath__63_0_I1795 (.Y(N5995), .A(N2579), .B(N6215));
NOR2XL inst_cellmath__63_0_I1796 (.Y(N6371), .A(N2579), .B(N5808));
NOR2XL inst_cellmath__63_0_I1797 (.Y(N5881), .A(N2579), .B(N6258));
NOR2XL inst_cellmath__63_0_I1798 (.Y(N6257), .A(N2579), .B(N5850));
NOR2XL inst_cellmath__63_0_I1799 (.Y(N5773), .A(N2579), .B(N6303));
NOR2XL inst_cellmath__63_0_I1800 (.Y(N6146), .A(N2579), .B(N5895));
NOR2XL inst_cellmath__63_0_I1801 (.Y(N6526), .A(N2579), .B(N6354));
NOR2XL inst_cellmath__63_0_I1802 (.Y(N6036), .A(N2579), .B(N5945));
NOR2XL inst_cellmath__63_0_I1803 (.Y(N6414), .A(N2579), .B(N6401));
NOR2XL inst_cellmath__63_0_I1804 (.Y(N5928), .A(N2579), .B(N5990));
NOR2XL inst_cellmath__63_0_I1805 (.Y(N6302), .A(N2579), .B(N6444));
NOR2XL inst_cellmath__63_0_I1806 (.Y(N5818), .A(N2579), .B(N6033));
NOR2XL inst_cellmath__63_0_I1808 (.Y(N5865), .A(N2648), .B(N6075));
NOR2XL inst_cellmath__63_0_I1809 (.Y(N6241), .A(N2648), .B(N6531));
NOR2XL inst_cellmath__63_0_I1810 (.Y(N5754), .A(N2648), .B(N6120));
NOR2XL inst_cellmath__63_0_I1811 (.Y(N6132), .A(N2648), .B(N6576));
NOR2XL inst_cellmath__63_0_I1812 (.Y(N6510), .A(N2648), .B(N6166));
NOR2XL inst_cellmath__63_0_I1813 (.Y(N6022), .A(N2648), .B(N5759));
NOR2XL inst_cellmath__63_0_I1814 (.Y(N6399), .A(N2648), .B(N6215));
NOR2XL inst_cellmath__63_0_I1815 (.Y(N5913), .A(N2648), .B(N5808));
NOR2XL inst_cellmath__63_0_I1816 (.Y(N6285), .A(N2648), .B(N6258));
NOR2XL inst_cellmath__63_0_I1817 (.Y(N5802), .A(N2648), .B(N5850));
NOR2XL inst_cellmath__63_0_I1818 (.Y(N6178), .A(N2648), .B(N6303));
NOR2XL inst_cellmath__63_0_I1819 (.Y(N6553), .A(N2648), .B(N5895));
NOR2XL inst_cellmath__63_0_I1820 (.Y(N6065), .A(N2648), .B(N6354));
NOR2XL inst_cellmath__63_0_I1821 (.Y(N6443), .A(N2648), .B(N5945));
NOR2XL inst_cellmath__63_0_I1822 (.Y(N5956), .A(N2648), .B(N6401));
NOR2XL inst_cellmath__63_0_I1823 (.Y(N6333), .A(N2648), .B(N5990));
NOR2XL inst_cellmath__63_0_I1824 (.Y(N5846), .A(N2648), .B(N6444));
NOR2XL inst_cellmath__63_0_I1825 (.Y(N6221), .A(N2648), .B(N6033));
NOR2XL inst_cellmath__63_0_I1827 (.Y(N6268), .A(N2746), .B(N6075));
NOR2XL inst_cellmath__63_0_I1828 (.Y(N5785), .A(N2746), .B(N6531));
NOR2XL inst_cellmath__63_0_I1829 (.Y(N6156), .A(N2746), .B(N6120));
NOR2XL inst_cellmath__63_0_I1830 (.Y(N6538), .A(N2746), .B(N6576));
NOR2XL inst_cellmath__63_0_I1831 (.Y(N6047), .A(N2746), .B(N6166));
NOR2XL inst_cellmath__63_0_I1832 (.Y(N6423), .A(N2746), .B(N5759));
NOR2XL inst_cellmath__63_0_I1833 (.Y(N5939), .A(N2746), .B(N6215));
NOR2XL inst_cellmath__63_0_I1834 (.Y(N6316), .A(N2746), .B(N5808));
NOR2XL inst_cellmath__63_0_I1835 (.Y(N5829), .A(N2746), .B(N6258));
NOR2XL inst_cellmath__63_0_I1836 (.Y(N6204), .A(N2746), .B(N5850));
NOR2XL inst_cellmath__63_0_I1837 (.Y(N5724), .A(N2746), .B(N6303));
NOR2XL inst_cellmath__63_0_I1838 (.Y(N6091), .A(N2746), .B(N5895));
NOR2XL inst_cellmath__63_0_I1839 (.Y(N6473), .A(N2746), .B(N6354));
NOR2XL inst_cellmath__63_0_I1840 (.Y(N5985), .A(N2746), .B(N5945));
NOR2XL inst_cellmath__63_0_I1841 (.Y(N6361), .A(N2746), .B(N6401));
NOR2XL inst_cellmath__63_0_I1842 (.Y(N5873), .A(N2746), .B(N5990));
NOR2XL inst_cellmath__63_0_I1843 (.Y(N6248), .A(N2746), .B(N6444));
NOR2XL inst_cellmath__63_0_I1844 (.Y(N5763), .A(N2746), .B(N6033));
NOR2XL inst_cellmath__63_0_I1846 (.Y(N5813), .A(N2822), .B(N6075));
NOR2XL inst_cellmath__63_0_I1847 (.Y(N6189), .A(N2822), .B(N6531));
NOR2XL inst_cellmath__63_0_I1848 (.Y(N6562), .A(N2822), .B(N6120));
NOR2XL inst_cellmath__63_0_I1849 (.Y(N6077), .A(N2822), .B(N6576));
NOR2XL inst_cellmath__63_0_I1850 (.Y(N6455), .A(N2822), .B(N6166));
NOR2XL inst_cellmath__63_0_I1851 (.Y(N5966), .A(N2822), .B(N5759));
NOR2XL inst_cellmath__63_0_I1852 (.Y(N6344), .A(N2822), .B(N6215));
NOR2XL inst_cellmath__63_0_I1853 (.Y(N5856), .A(N2822), .B(N5808));
NOR2XL inst_cellmath__63_0_I1854 (.Y(N6230), .A(N2822), .B(N6258));
NOR2XL inst_cellmath__63_0_I1855 (.Y(N5745), .A(N2822), .B(N5850));
NOR2XL inst_cellmath__63_0_I1856 (.Y(N6122), .A(N2822), .B(N6303));
NOR2XL inst_cellmath__63_0_I1857 (.Y(N6499), .A(N2822), .B(N5895));
NOR2XL inst_cellmath__63_0_I1858 (.Y(N6012), .A(N2822), .B(N6354));
NOR2XL inst_cellmath__63_0_I1859 (.Y(N6392), .A(N2822), .B(N5945));
NOR2XL inst_cellmath__63_0_I1860 (.Y(N5902), .A(N2822), .B(N6401));
NOR2XL inst_cellmath__63_0_I1861 (.Y(N6276), .A(N2822), .B(N5990));
NOR2XL inst_cellmath__63_0_I1862 (.Y(N5793), .A(N2822), .B(N6444));
NOR2XL inst_cellmath__63_0_I1863 (.Y(N6168), .A(N2822), .B(N6033));
NOR2XL inst_cellmath__63_0_I1865 (.Y(N6217), .A(N2887), .B(N6075));
NOR2XL inst_cellmath__63_0_I1866 (.Y(N5733), .A(N2887), .B(N6531));
NOR2XL inst_cellmath__63_0_I1867 (.Y(N6104), .A(N2887), .B(N6120));
NOR2XL inst_cellmath__63_0_I1868 (.Y(N6484), .A(N2887), .B(N6576));
NOR2XL inst_cellmath__63_0_I1869 (.Y(N5998), .A(N2887), .B(N6166));
NOR2XL inst_cellmath__63_0_I1870 (.Y(N6374), .A(N2887), .B(N5759));
NOR2XL inst_cellmath__63_0_I1871 (.Y(N5884), .A(N2887), .B(N6215));
NOR2XL inst_cellmath__63_0_I1872 (.Y(N6260), .A(N2887), .B(N5808));
NOR2XL inst_cellmath__63_0_I1873 (.Y(N5776), .A(N2887), .B(N6258));
NOR2XL inst_cellmath__63_0_I1874 (.Y(N6149), .A(N2887), .B(N5850));
NOR2XL inst_cellmath__63_0_I1875 (.Y(N6529), .A(N2887), .B(N6303));
NOR2XL inst_cellmath__63_0_I1876 (.Y(N6037), .A(N2887), .B(N5895));
NOR2XL inst_cellmath__63_0_I1877 (.Y(N6417), .A(N2887), .B(N6354));
NOR2XL inst_cellmath__63_0_I1878 (.Y(N5931), .A(N2887), .B(N5945));
NOR2XL inst_cellmath__63_0_I1879 (.Y(N6306), .A(N2887), .B(N6401));
NOR2XL inst_cellmath__63_0_I1880 (.Y(N5821), .A(N2887), .B(N5990));
NOR2XL inst_cellmath__63_0_I1881 (.Y(N6196), .A(N2887), .B(N6444));
NOR2XL inst_cellmath__63_0_I1882 (.Y(N6574), .A(N2887), .B(N6033));
NOR2XL inst_cellmath__63_0_I1884 (.Y(N5757), .A(N2637), .B(N6075));
NOR2XL inst_cellmath__63_0_I1885 (.Y(N6136), .A(N2637), .B(N6531));
NOR2XL inst_cellmath__63_0_I1886 (.Y(N6513), .A(N2637), .B(N6120));
NOR2XL inst_cellmath__63_0_I1887 (.Y(N6025), .A(N2637), .B(N6576));
NOR2XL inst_cellmath__63_0_I1888 (.Y(N6404), .A(N2637), .B(N6166));
NOR2XL inst_cellmath__63_0_I1889 (.Y(N5914), .A(N2637), .B(N5759));
NOR2XL inst_cellmath__63_0_I1890 (.Y(N6288), .A(N2637), .B(N6215));
NOR2XL inst_cellmath__63_0_I1891 (.Y(N5806), .A(N2637), .B(N5808));
NOR2XL inst_cellmath__63_0_I1892 (.Y(N6181), .A(N2637), .B(N6258));
NOR2XL inst_cellmath__63_0_I1893 (.Y(N6556), .A(N2637), .B(N5850));
NOR2XL inst_cellmath__63_0_I1894 (.Y(N6069), .A(N2637), .B(N6303));
NOR2XL inst_cellmath__63_0_I1895 (.Y(N6447), .A(N2637), .B(N5895));
NOR2XL inst_cellmath__63_0_I1896 (.Y(N5959), .A(N2637), .B(N6354));
NOR2XL inst_cellmath__63_0_I1897 (.Y(N6336), .A(N2637), .B(N5945));
NOR2XL inst_cellmath__63_0_I1898 (.Y(N5848), .A(N2637), .B(N6401));
NOR2XL inst_cellmath__63_0_I1899 (.Y(N6223), .A(N2637), .B(N5990));
NOR2XL inst_cellmath__63_0_I1900 (.Y(N5738), .A(N2637), .B(N6444));
NOR2XL inst_cellmath__63_0_I1901 (.Y(N6114), .A(N2637), .B(N6033));
NOR2XL inst_cellmath__63_0_I1903 (.Y(N6160), .A(N2705), .B(N6075));
NOR2XL inst_cellmath__63_0_I1904 (.Y(N6541), .A(N2705), .B(N6531));
NOR2XL inst_cellmath__63_0_I1905 (.Y(N6050), .A(N2705), .B(N6120));
NOR2XL inst_cellmath__63_0_I1906 (.Y(N6427), .A(N2705), .B(N6576));
NOR2XL inst_cellmath__63_0_I1907 (.Y(N5942), .A(N2705), .B(N6166));
NOR2XL inst_cellmath__63_0_I1908 (.Y(N6319), .A(N2705), .B(N5759));
NOR2XL inst_cellmath__63_0_I1909 (.Y(N5833), .A(N2705), .B(N6215));
NOR2XL inst_cellmath__63_0_I1910 (.Y(N6207), .A(N2705), .B(N5808));
NOR2XL inst_cellmath__63_0_I1911 (.Y(N5726), .A(N2705), .B(N6258));
NOR2XL inst_cellmath__63_0_I1912 (.Y(N6095), .A(N2705), .B(N5850));
NOR2XL inst_cellmath__63_0_I1913 (.Y(N6475), .A(N2705), .B(N6303));
NOR2XL inst_cellmath__63_0_I1914 (.Y(N5987), .A(N2705), .B(N5895));
NOR2XL inst_cellmath__63_0_I1915 (.Y(N6364), .A(N2705), .B(N6354));
NOR2XL inst_cellmath__63_0_I1916 (.Y(N5875), .A(N2705), .B(N5945));
NOR2XL inst_cellmath__63_0_I1917 (.Y(N6250), .A(N2705), .B(N6401));
NOR2XL inst_cellmath__63_0_I1918 (.Y(N5766), .A(N2705), .B(N5990));
NOR2XL inst_cellmath__63_0_I1919 (.Y(N6141), .A(N2705), .B(N6444));
NOR2XL inst_cellmath__63_0_I1920 (.Y(N6520), .A(N2705), .B(N6033));
NOR2XL inst_cellmath__63_0_I1922 (.Y(N6565), .A(N2776), .B(N6075));
NOR2XL inst_cellmath__63_0_I1923 (.Y(N6079), .A(N2776), .B(N6531));
NOR2XL inst_cellmath__63_0_I1924 (.Y(N6457), .A(N2776), .B(N6120));
NOR2XL inst_cellmath__63_0_I1925 (.Y(N5970), .A(N2776), .B(N6576));
NOR2XL inst_cellmath__63_0_I1926 (.Y(N6346), .A(N2776), .B(N6166));
NOR2XL inst_cellmath__63_0_I1927 (.Y(N5858), .A(N2776), .B(N5759));
NOR2XL inst_cellmath__63_0_I1928 (.Y(N6233), .A(N2776), .B(N6215));
NOR2XL inst_cellmath__63_0_I1929 (.Y(N5747), .A(N2776), .B(N5808));
NOR2XL inst_cellmath__63_0_I1930 (.Y(N6125), .A(N2776), .B(N6258));
NOR2XL inst_cellmath__63_0_I1931 (.Y(N6502), .A(N2776), .B(N5850));
NOR2XL inst_cellmath__63_0_I1932 (.Y(N6015), .A(N2776), .B(N6303));
NOR2XL inst_cellmath__63_0_I1933 (.Y(N6395), .A(N2776), .B(N5895));
NOR2XL inst_cellmath__63_0_I1934 (.Y(N5905), .A(N2776), .B(N6354));
NOR2XL inst_cellmath__63_0_I1935 (.Y(N6279), .A(N2776), .B(N5945));
NOR2XL inst_cellmath__63_0_I1936 (.Y(N5796), .A(N2776), .B(N6401));
NOR2XL inst_cellmath__63_0_I1937 (.Y(N6171), .A(N2776), .B(N5990));
NOR2XL inst_cellmath__63_0_I1938 (.Y(N6547), .A(N2776), .B(N6444));
NOR2XL inst_cellmath__63_0_I1939 (.Y(N6059), .A(N2776), .B(N6033));
NAND2XL inst_cellmath__63_0_I1940 (.Y(N6106), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[0]));
NAND2XL inst_cellmath__63_0_I1941 (.Y(N6486), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[1]));
NAND2XL inst_cellmath__63_0_I1942 (.Y(N6000), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[2]));
NAND2XL inst_cellmath__63_0_I1943 (.Y(N6376), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[3]));
NAND2XL inst_cellmath__63_0_I1944 (.Y(N5886), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[4]));
NAND2XL inst_cellmath__63_0_I1945 (.Y(N6262), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[5]));
NAND2XL inst_cellmath__63_0_I1946 (.Y(N5778), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[6]));
NAND2XL inst_cellmath__63_0_I1947 (.Y(N6151), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[7]));
NAND2XL inst_cellmath__63_0_I1948 (.Y(N6532), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[8]));
NAND2XL inst_cellmath__63_0_I1949 (.Y(N6039), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[9]));
NAND2XL inst_cellmath__63_0_I1950 (.Y(N6419), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[10]));
NAND2XL inst_cellmath__63_0_I1951 (.Y(N5932), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[11]));
NAND2XL inst_cellmath__63_0_I1952 (.Y(N6308), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[12]));
NAND2XL inst_cellmath__63_0_I1953 (.Y(N5823), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[13]));
NAND2XL inst_cellmath__63_0_I1954 (.Y(N6198), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[14]));
NAND2XL inst_cellmath__63_0_I1955 (.Y(N6577), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[15]));
NAND2XL inst_cellmath__63_0_I1956 (.Y(N6085), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[16]));
NAND2XL inst_cellmath__63_0_I1957 (.Y(N6466), .A(inst_cellmath__63__W0[33]), .B(inst_cellmath__51[17]));
ADDHX1 inst_cellmath__63_0_I1958 (.CO(N6102), .S(inst_cellmath__63__W1[2]), .A(N5969), .B(N6027));
ADDHX1 inst_cellmath__63_0_I1959 (.CO(N6483), .S(inst_cellmath__63__W0[3]), .A(N6377), .B(N6406));
ADDFX1 inst_cellmath__63_0_I1960 (.CO(N5996), .S(inst_cellmath__63__W1[3]), .A(N6430), .B(N6347), .CI(N6102));
ADDHX1 inst_cellmath__63_0_I1961 (.CO(N6372), .S(N6183), .A(N5916), .B(N5947));
ADDFX1 inst_cellmath__63_0_I1962 (.CO(N5882), .S(inst_cellmath__63__W0[4]), .A(N5859), .B(N5887), .CI(N5975));
ADDFX1 inst_cellmath__63_0_I1963 (.CO(inst_cellmath__63__W0[5]), .S(inst_cellmath__63__W1[4]), .A(N6183), .B(N6483), .CI(N5996));
ADDHX1 inst_cellmath__63_0_I1964 (.CO(N5774), .S(N6449), .A(N6232), .B(N6381));
ADDFX1 inst_cellmath__63_0_I1965 (.CO(N6147), .S(N5961), .A(N6263), .B(N6323), .CI(N6291));
ADDFX1 inst_cellmath__63_0_I1966 (.CO(N6527), .S(N6338), .A(N6372), .B(N6351), .CI(N6449));
ADDFX1 inst_cellmath__63_0_I1967 (.CO(inst_cellmath__63__W0[6]), .S(inst_cellmath__63__W1[5]), .A(N5961), .B(N5882), .CI(N6338));
ADDHX1 inst_cellmath__63_0_I1968 (.CO(N6415), .S(N6226), .A(N5779), .B(N5919));
ADDFX1 inst_cellmath__63_0_I1969 (.CO(N5929), .S(N5740), .A(N5809), .B(N5863), .CI(N5836));
ADDFX1 inst_cellmath__63_0_I1970 (.CO(N6304), .S(N6115), .A(N5890), .B(N5748), .CI(N5774));
ADDFX1 inst_cellmath__63_0_I1971 (.CO(N5819), .S(N6493), .A(N6226), .B(N6147), .CI(N5740));
ADDFX1 inst_cellmath__63_0_I1972 (.CO(inst_cellmath__63__W0[7]), .S(inst_cellmath__63__W1[6]), .A(N6115), .B(N6527), .CI(N6493));
ADDHX1 inst_cellmath__63_0_I1973 (.CO(N6572), .S(N6386), .A(N6184), .B(N6326));
ADDFX1 inst_cellmath__63_0_I1974 (.CO(N6083), .S(N5896), .A(N6211), .B(N6266), .CI(N6126));
ADDFX1 inst_cellmath__63_0_I1975 (.CO(N6462), .S(N6271), .A(N6152), .B(N6238), .CI(N6293));
ADDFX1 inst_cellmath__63_0_I1976 (.CO(N5977), .S(N5789), .A(N5929), .B(N6415), .CI(N6386));
ADDFX1 inst_cellmath__63_0_I1977 (.CO(N6355), .S(N6162), .A(N6304), .B(N5896), .CI(N6271));
ADDFX1 inst_cellmath__63_0_I1978 (.CO(inst_cellmath__63__W0[8]), .S(inst_cellmath__63__W1[7]), .A(N5789), .B(N5819), .CI(N6162));
ADDHX1 inst_cellmath__63_0_I1979 (.CO(N6242), .S(N6053), .A(N5728), .B(N5865));
ADDFX1 inst_cellmath__63_0_I1980 (.CO(N5756), .S(N6431), .A(N5752), .B(N5811), .CI(N6501));
ADDFX1 inst_cellmath__63_0_I1981 (.CO(N6134), .S(N5946), .A(N6533), .B(N5783), .CI(N6558));
ADDFX1 inst_cellmath__63_0_I1982 (.CO(N6511), .S(N6322), .A(N6572), .B(N5839), .CI(N6053));
ADDFX1 inst_cellmath__63_0_I1983 (.CO(N6024), .S(N5837), .A(N6462), .B(N6083), .CI(N6431));
ADDFX1 inst_cellmath__63_0_I1984 (.CO(N6402), .S(N6210), .A(N5977), .B(N5946), .CI(N6322));
ADDFX1 inst_cellmath__63_0_I1985 (.CO(inst_cellmath__63__W0[9]), .S(inst_cellmath__63__W1[8]), .A(N5837), .B(N6355), .CI(N6210));
ADDHX1 inst_cellmath__63_0_I1986 (.CO(N6287), .S(N6099), .A(N6130), .B(N6268));
ADDFX1 inst_cellmath__63_0_I1987 (.CO(N5804), .S(N6478), .A(N6016), .B(N6214), .CI(N6040));
ADDFX1 inst_cellmath__63_0_I1988 (.CO(N6179), .S(N5991), .A(N6155), .B(N6187), .CI(N6071));
ADDFX1 inst_cellmath__63_0_I1989 (.CO(N6555), .S(N6368), .A(N6241), .B(N6098), .CI(N6242));
ADDFX1 inst_cellmath__63_0_I1990 (.CO(N6067), .S(N5878), .A(N5756), .B(N6099), .CI(N6134));
ADDFX1 inst_cellmath__63_0_I1991 (.CO(N6445), .S(N6253), .A(N6478), .B(N5991), .CI(N6511));
ADDFX1 inst_cellmath__63_0_I1992 (.CO(N5958), .S(N5770), .A(N6024), .B(N6368), .CI(N5878));
ADDFX1 inst_cellmath__63_0_I1993 (.CO(inst_cellmath__63__W0[10]), .S(inst_cellmath__63__W1[9]), .A(N6253), .B(N6402), .CI(N5770));
ADDHX1 inst_cellmath__63_0_I1994 (.CO(N5847), .S(N6522), .A(N6536), .B(N5813));
ADDFX1 inst_cellmath__63_0_I1995 (.CO(N6222), .S(N6034), .A(N6420), .B(N5754), .CI(N6450));
ADDFX1 inst_cellmath__63_0_I1996 (.CO(N5737), .S(N6411), .A(N6560), .B(N6396), .CI(N6479));
ADDFX1 inst_cellmath__63_0_I1997 (.CO(N6113), .S(N5926), .A(N6507), .B(N5731), .CI(N5785));
ADDFX1 inst_cellmath__63_0_I1998 (.CO(N6490), .S(N6300), .A(N6522), .B(N6287), .CI(N5804));
ADDFX1 inst_cellmath__63_0_I1999 (.CO(N6005), .S(N5816), .A(N6411), .B(N6179), .CI(N6034));
ADDFX1 inst_cellmath__63_0_I2000 (.CO(N6384), .S(N6193), .A(N5926), .B(N6555), .CI(N6067));
ADDFX1 inst_cellmath__63_0_I2001 (.CO(N5893), .S(N6569), .A(N6445), .B(N6300), .CI(N5816));
ADDFX1 inst_cellmath__63_0_I2002 (.CO(inst_cellmath__63__W0[11]), .S(inst_cellmath__63__W1[10]), .A(N5958), .B(N6193), .CI(N6569));
ADDHX1 inst_cellmath__63_0_I2003 (.CO(N5787), .S(N6460), .A(N6074), .B(N6217));
ADDFX1 inst_cellmath__63_0_I2004 (.CO(N6159), .S(N5974), .A(N5962), .B(N6156), .CI(N5992));
ADDFX1 inst_cellmath__63_0_I2005 (.CO(N6540), .S(N6350), .A(N6101), .B(N5933), .CI(N6020));
ADDFX1 inst_cellmath__63_0_I2006 (.CO(N6049), .S(N5862), .A(N6045), .B(N6132), .CI(N6189));
ADDFX1 inst_cellmath__63_0_I2007 (.CO(N6426), .S(N6237), .A(N5847), .B(N5904), .CI(N6460));
ADDFX1 inst_cellmath__63_0_I2008 (.CO(N5941), .S(N5751), .A(N6222), .B(N5737), .CI(N6113));
ADDFX1 inst_cellmath__63_0_I2009 (.CO(N6318), .S(N6129), .A(N5974), .B(N6350), .CI(N5862));
ADDFX1 inst_cellmath__63_0_I2010 (.CO(N5832), .S(N6506), .A(N6237), .B(N6490), .CI(N6005));
ADDFX1 inst_cellmath__63_0_I2011 (.CO(N6206), .S(N6019), .A(N6384), .B(N5751), .CI(N6129));
ADDFX1 inst_cellmath__63_0_I2012 (.CO(inst_cellmath__63__W0[12]), .S(inst_cellmath__63__W1[11]), .A(N5893), .B(N6506), .CI(N6019));
ADDHX1 inst_cellmath__63_0_I2013 (.CO(N6094), .S(N5909), .A(N6482), .B(N5757));
ADDFX1 inst_cellmath__63_0_I2014 (.CO(N6474), .S(N6282), .A(N6367), .B(N6562), .CI(N6398));
ADDFX1 inst_cellmath__63_0_I2015 (.CO(N5986), .S(N5799), .A(N6510), .B(N6339), .CI(N6422));
ADDFX1 inst_cellmath__63_0_I2016 (.CO(N6363), .S(N6174), .A(N6453), .B(N6538), .CI(N6309));
ADDFX1 inst_cellmath__63_0_I2017 (.CO(N5874), .S(N6550), .A(N5733), .B(N6280), .CI(N5787));
ADDFX1 inst_cellmath__63_0_I2018 (.CO(N6249), .S(N6062), .A(N6540), .B(N5909), .CI(N6159));
ADDFX1 inst_cellmath__63_0_I2019 (.CO(N5765), .S(N6439), .A(N5799), .B(N6049), .CI(N6282));
ADDFX1 inst_cellmath__63_0_I2020 (.CO(N6140), .S(N5953), .A(N6426), .B(N6174), .CI(N5941));
ADDFX1 inst_cellmath__63_0_I2021 (.CO(N6519), .S(N6330), .A(N6062), .B(N6550), .CI(N6318));
ADDFX1 inst_cellmath__63_0_I2022 (.CO(N6030), .S(N5844), .A(N5832), .B(N6439), .CI(N5953));
ADDFX1 inst_cellmath__63_0_I2023 (.CO(inst_cellmath__63__W0[13]), .S(inst_cellmath__63__W1[12]), .A(N6330), .B(N6206), .CI(N5844));
ADDHX1 inst_cellmath__63_0_I2024 (.CO(N5922), .S(N5735), .A(N6022), .B(N6160));
ADDFX1 inst_cellmath__63_0_I2025 (.CO(N6296), .S(N6109), .A(N5797), .B(N6104), .CI(N5937));
ADDFX1 inst_cellmath__63_0_I2026 (.CO(N5814), .S(N6488), .A(N5910), .B(N5879), .CI(N5964));
ADDFX1 inst_cellmath__63_0_I2027 (.CO(N6190), .S(N6002), .A(N6047), .B(N6077), .CI(N5995));
ADDFX1 inst_cellmath__63_0_I2028 (.CO(N6564), .S(N6380), .A(N6136), .B(N5824), .CI(N5851));
ADDFX1 inst_cellmath__63_0_I2029 (.CO(N6078), .S(N5889), .A(N5735), .B(N6094), .CI(N6474));
ADDFX1 inst_cellmath__63_0_I2030 (.CO(N6456), .S(N6265), .A(N6363), .B(N5986), .CI(N6488));
ADDFX1 inst_cellmath__63_0_I2031 (.CO(N5968), .S(N5782), .A(N6002), .B(N6109), .CI(N5874));
ADDFX1 inst_cellmath__63_0_I2032 (.CO(N6345), .S(N6154), .A(N6249), .B(N6380), .CI(N5765));
ADDFX1 inst_cellmath__63_0_I2033 (.CO(N5857), .S(N6535), .A(N6265), .B(N5889), .CI(N6140));
ADDFX1 inst_cellmath__63_0_I2034 (.CO(N6231), .S(N6044), .A(N6519), .B(N5782), .CI(N6154));
ADDFX1 inst_cellmath__63_0_I2035 (.CO(inst_cellmath__63__W0[14]), .S(inst_cellmath__63__W1[13]), .A(N6030), .B(N6535), .CI(N6044));
ADDHX1 inst_cellmath__63_0_I2036 (.CO(N6124), .S(N5936), .A(N6170), .B(N6199));
ADDFX1 inst_cellmath__63_0_I2037 (.CO(N6500), .S(N6313), .A(N6513), .B(N6423), .CI(N6342));
ADDFX1 inst_cellmath__63_0_I2038 (.CO(N6014), .S(N5827), .A(N6314), .B(N6283), .CI(N6371));
ADDFX1 inst_cellmath__63_0_I2039 (.CO(N6394), .S(N6202), .A(N6455), .B(N6484), .CI(N6399));
ADDFX1 inst_cellmath__63_0_I2040 (.CO(N5903), .S(N5721), .A(N6565), .B(N6225), .CI(N6254));
ADDFX1 inst_cellmath__63_0_I2041 (.CO(N6278), .S(N6089), .A(N5922), .B(N6541), .CI(N5936));
ADDFX1 inst_cellmath__63_0_I2042 (.CO(N5795), .S(N6470), .A(N6190), .B(N5814), .CI(N6296));
ADDFX1 inst_cellmath__63_0_I2043 (.CO(N6169), .S(N5982), .A(N5827), .B(N6564), .CI(N6202));
ADDFX1 inst_cellmath__63_0_I2044 (.CO(N6546), .S(N6360), .A(N5721), .B(N6313), .CI(N6078));
ADDFX1 inst_cellmath__63_0_I2045 (.CO(N6058), .S(N5870), .A(N6456), .B(N6089), .CI(N6470));
ADDFX1 inst_cellmath__63_0_I2046 (.CO(N6435), .S(N6246), .A(N5982), .B(N5968), .CI(N6360));
ADDFX1 inst_cellmath__63_0_I2047 (.CO(N5950), .S(N5762), .A(N5870), .B(N6345), .CI(N5857));
ADDFX1 inst_cellmath__63_0_I2048 (.CO(inst_cellmath__63__W0[15]), .S(inst_cellmath__63__W1[14]), .A(N6246), .B(N6231), .CI(N5762));
XNOR2X1 inst_cellmath__63_0_I2049 (.Y(N6516), .A(N6106), .B(N6548));
OR2XL inst_cellmath__63_0_I2050 (.Y(N5841), .A(N6106), .B(N6548));
ADDFX1 inst_cellmath__63_0_I2051 (.CO(N5734), .S(N6408), .A(N5966), .B(N6578), .CI(N5881));
ADDFX1 inst_cellmath__63_0_I2052 (.CO(N6105), .S(N5918), .A(N5741), .B(N6050), .CI(N5913));
ADDFX1 inst_cellmath__63_0_I2053 (.CO(N6485), .S(N6294), .A(N5854), .B(N5828), .CI(N5998));
ADDFX1 inst_cellmath__63_0_I2054 (.CO(N5999), .S(N5810), .A(N5939), .B(N6025), .CI(N5800));
ADDFX1 inst_cellmath__63_0_I2055 (.CO(N6375), .S(N6186), .A(N6079), .B(N5769), .CI(N6124));
ADDFX1 inst_cellmath__63_0_I2056 (.CO(N5885), .S(N6561), .A(N6014), .B(N6516), .CI(N6394));
ADDFX1 inst_cellmath__63_0_I2057 (.CO(N6261), .S(N6073), .A(N5903), .B(N6500), .CI(N6294));
ADDFX1 inst_cellmath__63_0_I2058 (.CO(N5777), .S(N6452), .A(N6408), .B(N5918), .CI(N5810));
ADDFX1 inst_cellmath__63_0_I2059 (.CO(N6150), .S(N5965), .A(N6186), .B(N6278), .CI(N5795));
ADDFX1 inst_cellmath__63_0_I2060 (.CO(N6530), .S(N6341), .A(N6169), .B(N6561), .CI(N6073));
ADDFX1 inst_cellmath__63_0_I2061 (.CO(N6038), .S(N5853), .A(N6452), .B(N6546), .CI(N6058));
ADDFX1 inst_cellmath__63_0_I2062 (.CO(N6418), .S(N6228), .A(N6341), .B(N5965), .CI(N6435));
ADDFX1 inst_cellmath__63_0_I2063 (.CO(inst_cellmath__63__W0[16]), .S(inst_cellmath__63__W1[15]), .A(N5950), .B(N5853), .CI(N6228));
ADDFX1 inst_cellmath__63_0_I2064 (.CO(N6307), .S(N6118), .A(N6486), .B(N6060), .CI(N6086));
ADDFX1 inst_cellmath__63_0_I2065 (.CO(N5822), .S(N6496), .A(N6374), .B(N6116), .CI(N6285));
ADDFX1 inst_cellmath__63_0_I2066 (.CO(N6197), .S(N6009), .A(N6144), .B(N6457), .CI(N6316));
ADDFX1 inst_cellmath__63_0_I2067 (.CO(N6575), .S(N6389), .A(N6257), .B(N6227), .CI(N6404));
ADDFX1 inst_cellmath__63_0_I2068 (.CO(N6084), .S(N5899), .A(N6344), .B(N6427), .CI(N6203));
ADDFX1 inst_cellmath__63_0_I2069 (.CO(N6465), .S(N6273), .A(N5841), .B(N6175), .CI(N6485));
ADDFX1 inst_cellmath__63_0_I2070 (.CO(N5979), .S(N5791), .A(N5734), .B(N6105), .CI(N6118));
ADDFX1 inst_cellmath__63_0_I2071 (.CO(N6357), .S(N6165), .A(N6375), .B(N5999), .CI(N6496));
ADDFX1 inst_cellmath__63_0_I2072 (.CO(N5868), .S(N6545), .A(N6009), .B(N6389), .CI(N5899));
ADDFX1 inst_cellmath__63_0_I2073 (.CO(N6244), .S(N6055), .A(N6261), .B(N5885), .CI(N6273));
ADDFX1 inst_cellmath__63_0_I2074 (.CO(N5758), .S(N6433), .A(N5777), .B(N5791), .CI(N6165));
ADDFX1 inst_cellmath__63_0_I2075 (.CO(N6137), .S(N5948), .A(N6545), .B(N6150), .CI(N6530));
ADDFX1 inst_cellmath__63_0_I2076 (.CO(N6514), .S(N6325), .A(N6038), .B(N6055), .CI(N6433));
ADDFX1 inst_cellmath__63_0_I2077 (.CO(inst_cellmath__63__W0[17]), .S(inst_cellmath__63__W1[16]), .A(N6418), .B(N5948), .CI(N6325));
ADDFX1 inst_cellmath__63_0_I2078 (.CO(N6405), .S(N6213), .A(N6000), .B(N6436), .CI(N6467));
ADDFX1 inst_cellmath__63_0_I2079 (.CO(N5915), .S(N5730), .A(N6523), .B(N6492), .CI(N5914));
ADDFX1 inst_cellmath__63_0_I2080 (.CO(N6290), .S(N6100), .A(N6551), .B(N5773), .CI(N5829));
ADDFX1 inst_cellmath__63_0_I2081 (.CO(N5807), .S(N6481), .A(N5802), .B(N5970), .CI(N5856));
ADDFX1 inst_cellmath__63_0_I2082 (.CO(N6182), .S(N5994), .A(N5884), .B(N5942), .CI(N5743));
ADDFX1 inst_cellmath__63_0_I2083 (.CO(N6557), .S(N6370), .A(N6213), .B(N5722), .CI(N6307));
ADDFX1 inst_cellmath__63_0_I2084 (.CO(N6070), .S(N5880), .A(N6197), .B(N6575), .CI(N5822));
ADDFX1 inst_cellmath__63_0_I2085 (.CO(N6448), .S(N6256), .A(N5730), .B(N6084), .CI(N6481));
ADDFX1 inst_cellmath__63_0_I2086 (.CO(N5960), .S(N5772), .A(N5994), .B(N6100), .CI(N6465));
ADDFX1 inst_cellmath__63_0_I2087 (.CO(N6337), .S(N6145), .A(N6370), .B(N5979), .CI(N6357));
ADDFX1 inst_cellmath__63_0_I2088 (.CO(N5849), .S(N6525), .A(N5868), .B(N5880), .CI(N6256));
ADDFX1 inst_cellmath__63_0_I2089 (.CO(N6224), .S(N6035), .A(N6244), .B(N5772), .CI(N6145));
ADDFX1 inst_cellmath__63_0_I2090 (.CO(N5739), .S(N6413), .A(N6525), .B(N5758), .CI(N6137));
ADDFX1 inst_cellmath__63_0_I2091 (.CO(inst_cellmath__63__W0[18]), .S(inst_cellmath__63__W1[17]), .A(N6514), .B(N6035), .CI(N6413));
INVXL inst_cellmath__63_0_I2092 (.Y(N5920), .A(N6299));
ADDFX1 inst_cellmath__63_0_I2093 (.CO(N6491), .S(N6301), .A(N6376), .B(N5980), .CI(N5920));
ADDFX1 inst_cellmath__63_0_I2094 (.CO(N6385), .S(N6194), .A(N6032), .B(N6007), .CI(N6063));
ADDFX1 inst_cellmath__63_0_I2095 (.CO(N5894), .S(N6570), .A(N6178), .B(N6319), .CI(N6230));
ADDFX1 inst_cellmath__63_0_I2096 (.CO(N6270), .S(N6082), .A(N6090), .B(N6346), .CI(N6119));
ADDFX1 inst_cellmath__63_0_I2097 (.CO(N5788), .S(N6461), .A(N6260), .B(N6204), .CI(N6288));
ADDFX1 inst_cellmath__63_0_I2098 (.CO(N6161), .S(N5976), .A(N6146), .B(N6405), .CI(N6301));
ADDFX1 inst_cellmath__63_0_I2099 (.CO(N6543), .S(N6352), .A(N5807), .B(N5915), .CI(N6290));
ADDFX1 inst_cellmath__63_0_I2100 (.CO(N6051), .S(N5864), .A(N6182), .B(N6194), .CI(N6570));
ADDFX1 inst_cellmath__63_0_I2101 (.CO(N6428), .S(N6240), .A(N6082), .B(N6461), .CI(N6557));
ADDFX1 inst_cellmath__63_0_I2102 (.CO(N5944), .S(N5753), .A(N5976), .B(N6070), .CI(N6448));
ADDFX1 inst_cellmath__63_0_I2103 (.CO(N6320), .S(N6131), .A(N5960), .B(N6352), .CI(N5864));
ADDFX1 inst_cellmath__63_0_I2104 (.CO(N5834), .S(N6509), .A(N6337), .B(N6240), .CI(N5753));
ADDFX1 inst_cellmath__63_0_I2105 (.CO(N6209), .S(N6021), .A(N6131), .B(N5849), .CI(N6224));
ADDFX1 inst_cellmath__63_0_I2106 (.CO(inst_cellmath__63__W0[19]), .S(inst_cellmath__63__W1[18]), .A(N5739), .B(N6509), .CI(N6021));
ADDFX1 inst_cellmath__63_0_I2107 (.CO(N6096), .S(N5912), .A(N6299), .B(N6568), .CI(N6387));
ADDFX1 inst_cellmath__63_0_I2108 (.CO(N6477), .S(N6284), .A(N6412), .B(N5886), .CI(N5912));
ADDFX1 inst_cellmath__63_0_I2109 (.CO(N5988), .S(N5801), .A(N6471), .B(N6440), .CI(N5858));
ADDFX1 inst_cellmath__63_0_I2110 (.CO(N6365), .S(N6177), .A(N6491), .B(N5724), .CI(N5776));
ADDFX1 inst_cellmath__63_0_I2111 (.CO(N5877), .S(N6552), .A(N6495), .B(N5745), .CI(N6526));
ADDFX1 inst_cellmath__63_0_I2112 (.CO(N6251), .S(N6064), .A(N5833), .B(N5806), .CI(N6553));
ADDFX1 inst_cellmath__63_0_I2113 (.CO(N5767), .S(N6442), .A(N6284), .B(N6385), .CI(N5894));
ADDFX1 inst_cellmath__63_0_I2114 (.CO(N6143), .S(N5955), .A(N6270), .B(N5788), .CI(N5801));
ADDFX1 inst_cellmath__63_0_I2115 (.CO(N6521), .S(N6332), .A(N6161), .B(N6552), .CI(N6064));
ADDFX1 inst_cellmath__63_0_I2116 (.CO(N6031), .S(N5845), .A(N6543), .B(N6177), .CI(N6051));
ADDFX1 inst_cellmath__63_0_I2117 (.CO(N6410), .S(N6220), .A(N6428), .B(N6442), .CI(N5955));
ADDFX1 inst_cellmath__63_0_I2118 (.CO(N5925), .S(N5736), .A(N5944), .B(N6332), .CI(N5845));
ADDFX1 inst_cellmath__63_0_I2119 (.CO(N6297), .S(N6110), .A(N6220), .B(N6320), .CI(N5834));
ADDFX1 inst_cellmath__63_0_I2120 (.CO(inst_cellmath__63__W0[20]), .S(inst_cellmath__63__W1[19]), .A(N6209), .B(N5736), .CI(N6110));
ADDFX1 inst_cellmath__63_0_I2121 (.CO(N6192), .S(N6003), .A(N5927), .B(N5973), .CI(N6096));
ADDFX1 inst_cellmath__63_0_I2122 (.CO(N6566), .S(N6382), .A(N5954), .B(N6262), .CI(N5983));
ADDFX1 inst_cellmath__63_0_I2123 (.CO(N6080), .S(N5892), .A(N6122), .B(N6010), .CI(N6181));
ADDFX1 inst_cellmath__63_0_I2124 (.CO(N6459), .S(N6267), .A(N6036), .B(N6149), .CI(N6065));
ADDFX1 inst_cellmath__63_0_I2125 (.CO(N5971), .S(N5784), .A(N6233), .B(N6207), .CI(N6091));
ADDFX1 inst_cellmath__63_0_I2126 (.CO(N6348), .S(N6158), .A(N6003), .B(N6477), .CI(N5988));
ADDFX1 inst_cellmath__63_0_I2127 (.CO(N5861), .S(N6537), .A(N6382), .B(N5877), .CI(N6251));
ADDFX1 inst_cellmath__63_0_I2128 (.CO(N6234), .S(N6046), .A(N5892), .B(N6365), .CI(N6267));
ADDFX1 inst_cellmath__63_0_I2129 (.CO(N5749), .S(N6425), .A(N5767), .B(N5784), .CI(N6143));
ADDFX1 inst_cellmath__63_0_I2130 (.CO(N6128), .S(N5938), .A(N6521), .B(N6158), .CI(N6537));
ADDFX1 inst_cellmath__63_0_I2131 (.CO(N6503), .S(N6315), .A(N6031), .B(N6046), .CI(N6425));
ADDFX1 inst_cellmath__63_0_I2132 (.CO(N6017), .S(N5831), .A(N5938), .B(N6410), .CI(N5925));
ADDFX1 inst_cellmath__63_0_I2133 (.CO(inst_cellmath__63__W0[21]), .S(inst_cellmath__63__W1[20]), .A(N6297), .B(N6315), .CI(N5831));
ADDFX1 inst_cellmath__63_0_I2134 (.CO(N5906), .S(N5723), .A(N6331), .B(N2875), .CI(N5778));
ADDFX1 inst_cellmath__63_0_I2135 (.CO(N6281), .S(N6093), .A(N6390), .B(N6359), .CI(N6414));
ADDFX1 inst_cellmath__63_0_I2136 (.CO(N5798), .S(N6472), .A(N6529), .B(N6192), .CI(N5726));
ADDFX1 inst_cellmath__63_0_I2137 (.CO(N6172), .S(N5984), .A(N6443), .B(N6556), .CI(N6473));
ADDFX1 inst_cellmath__63_0_I2138 (.CO(N6549), .S(N6362), .A(N6499), .B(N5747), .CI(N5723));
ADDFX1 inst_cellmath__63_0_I2139 (.CO(N6061), .S(N5872), .A(N6080), .B(N6566), .CI(N6459));
ADDFX1 inst_cellmath__63_0_I2140 (.CO(N6437), .S(N6247), .A(N5971), .B(N6093), .CI(N6472));
ADDFX1 inst_cellmath__63_0_I2141 (.CO(N5952), .S(N5764), .A(N6348), .B(N5984), .CI(N6362));
ADDFX1 inst_cellmath__63_0_I2142 (.CO(N6329), .S(N6139), .A(N5872), .B(N5861), .CI(N6234));
ADDFX1 inst_cellmath__63_0_I2143 (.CO(N5842), .S(N6517), .A(N5749), .B(N6247), .CI(N5764));
ADDFX1 inst_cellmath__63_0_I2144 (.CO(N6218), .S(N6029), .A(N6139), .B(N6128), .CI(N6503));
ADDFX1 inst_cellmath__63_0_I2145 (.CO(inst_cellmath__63__W0[22]), .S(inst_cellmath__63__W1[21]), .A(N6017), .B(N6517), .CI(N6029));
ADDFX1 inst_cellmath__63_0_I2146 (.CO(N6107), .S(N5921), .A(N5871), .B(N2631), .CI(N6151));
ADDFX1 inst_cellmath__63_0_I2147 (.CO(N6487), .S(N6295), .A(N5928), .B(N5898), .CI(N5956));
ADDFX1 inst_cellmath__63_0_I2148 (.CO(N6001), .S(N5812), .A(N5906), .B(N6069), .CI(N6125));
ADDFX1 inst_cellmath__63_0_I2149 (.CO(N6378), .S(N6188), .A(N5985), .B(N6095), .CI(N6012));
ADDFX1 inst_cellmath__63_0_I2150 (.CO(N5888), .S(N6563), .A(N5921), .B(N6037), .CI(N6281));
ADDFX1 inst_cellmath__63_0_I2151 (.CO(N6264), .S(N6076), .A(N6172), .B(N5798), .CI(N6295));
ADDFX1 inst_cellmath__63_0_I2152 (.CO(N5780), .S(N6454), .A(N6188), .B(N6549), .CI(N5812));
ADDFX1 inst_cellmath__63_0_I2153 (.CO(N6153), .S(N5967), .A(N6563), .B(N6061), .CI(N6437));
ADDFX1 inst_cellmath__63_0_I2154 (.CO(N6534), .S(N6343), .A(N5952), .B(N6076), .CI(N6454));
ADDFX1 inst_cellmath__63_0_I2155 (.CO(N6041), .S(N5855), .A(N5967), .B(N6329), .CI(N5842));
ADDFX1 inst_cellmath__63_0_I2156 (.CO(inst_cellmath__63__W0[23]), .S(inst_cellmath__63__W1[22]), .A(N6218), .B(N6343), .CI(N5855));
ADDFX1 inst_cellmath__63_0_I2157 (.CO(N5935), .S(N5744), .A(N6274), .B(N2698), .CI(N6532));
ADDFX1 inst_cellmath__63_0_I2158 (.CO(N6310), .S(N6121), .A(N6333), .B(N6302), .CI(N6361));
ADDFX1 inst_cellmath__63_0_I2159 (.CO(N5825), .S(N6498), .A(N6475), .B(N6107), .CI(N6392));
ADDFX1 inst_cellmath__63_0_I2160 (.CO(N6201), .S(N6011), .A(N6417), .B(N6502), .CI(N6447));
ADDFX1 inst_cellmath__63_0_I2161 (.CO(N6579), .S(N6391), .A(N6487), .B(N5744), .CI(N6378));
ADDFX1 inst_cellmath__63_0_I2162 (.CO(N6087), .S(N5901), .A(N6121), .B(N6001), .CI(N6498));
ADDFX1 inst_cellmath__63_0_I2163 (.CO(N6469), .S(N6275), .A(N6011), .B(N5888), .CI(N6264));
ADDFX1 inst_cellmath__63_0_I2164 (.CO(N5981), .S(N5792), .A(N5780), .B(N6391), .CI(N5901));
ADDFX1 inst_cellmath__63_0_I2165 (.CO(N6358), .S(N6167), .A(N6275), .B(N6153), .CI(N6534));
ADDFX1 inst_cellmath__63_0_I2166 (.CO(inst_cellmath__63__W0[24]), .S(inst_cellmath__63__W1[23]), .A(N6041), .B(N5792), .CI(N6167));
ADDFX1 inst_cellmath__63_0_I2167 (.CO(N6245), .S(N6056), .A(N5818), .B(N2772), .CI(N6039));
ADDFX1 inst_cellmath__63_0_I2168 (.CO(N5760), .S(N6434), .A(N5873), .B(N5846), .CI(N5902));
ADDFX1 inst_cellmath__63_0_I2169 (.CO(N6138), .S(N5949), .A(N6015), .B(N5935), .CI(N5931));
ADDFX1 inst_cellmath__63_0_I2170 (.CO(N6515), .S(N6327), .A(N5987), .B(N5959), .CI(N6056));
ADDFX1 inst_cellmath__63_0_I2171 (.CO(N6028), .S(N5840), .A(N5825), .B(N6310), .CI(N6434));
ADDFX1 inst_cellmath__63_0_I2172 (.CO(N6407), .S(N6216), .A(N5949), .B(N6201), .CI(N6327));
ADDFX1 inst_cellmath__63_0_I2173 (.CO(N5917), .S(N5732), .A(N6087), .B(N6579), .CI(N5840));
ADDFX1 inst_cellmath__63_0_I2174 (.CO(N6292), .S(N6103), .A(N6216), .B(N6469), .CI(N5981));
ADDFX1 inst_cellmath__63_0_I2175 (.CO(inst_cellmath__63__W0[25]), .S(inst_cellmath__63__W1[24]), .A(N6358), .B(N5732), .CI(N6103));
ADDFX1 inst_cellmath__63_0_I2176 (.CO(N6185), .S(N5997), .A(N6221), .B(N2579), .CI(N6419));
ADDFX1 inst_cellmath__63_0_I2177 (.CO(N6559), .S(N6373), .A(N6276), .B(N6248), .CI(N6306));
ADDFX1 inst_cellmath__63_0_I2178 (.CO(N6072), .S(N5883), .A(N6336), .B(N6245), .CI(N6364));
ADDFX1 inst_cellmath__63_0_I2179 (.CO(N6451), .S(N6259), .A(N5997), .B(N6395), .CI(N5760));
ADDFX1 inst_cellmath__63_0_I2180 (.CO(N5963), .S(N5775), .A(N6373), .B(N6138), .CI(N6515));
ADDFX1 inst_cellmath__63_0_I2181 (.CO(N6340), .S(N6148), .A(N6259), .B(N5883), .CI(N6028));
ADDFX1 inst_cellmath__63_0_I2182 (.CO(N5852), .S(N6528), .A(N6407), .B(N5775), .CI(N5917));
ADDFX1 inst_cellmath__63_0_I2183 (.CO(inst_cellmath__63__W0[26]), .S(inst_cellmath__63__W1[25]), .A(N6292), .B(N6148), .CI(N6528));
ADDFX1 inst_cellmath__63_0_I2184 (.CO(N5742), .S(N6416), .A(N5763), .B(N2648), .CI(N5793));
ADDFX1 inst_cellmath__63_0_I2185 (.CO(N6117), .S(N5930), .A(N5821), .B(N5932), .CI(N5848));
ADDFX1 inst_cellmath__63_0_I2186 (.CO(N6494), .S(N6305), .A(N5875), .B(N6185), .CI(N5905));
ADDFX1 inst_cellmath__63_0_I2187 (.CO(N6008), .S(N5820), .A(N6559), .B(N6416), .CI(N6072));
ADDFX1 inst_cellmath__63_0_I2188 (.CO(N6388), .S(N6195), .A(N6305), .B(N5930), .CI(N6451));
ADDFX1 inst_cellmath__63_0_I2189 (.CO(N5897), .S(N6573), .A(N5820), .B(N5963), .CI(N6195));
ADDFX1 inst_cellmath__63_0_I2190 (.CO(inst_cellmath__63__W1[27]), .S(inst_cellmath__63__W1[26]), .A(N5852), .B(N6340), .CI(N6573));
ADDFX1 inst_cellmath__63_0_I2191 (.CO(N5790), .S(N6463), .A(N6168), .B(N2746), .CI(N6308));
ADDFX1 inst_cellmath__63_0_I2192 (.CO(N6163), .S(N5978), .A(N6223), .B(N6196), .CI(N6250));
ADDFX1 inst_cellmath__63_0_I2193 (.CO(N6544), .S(N6356), .A(N5742), .B(N6279), .CI(N6463));
ADDFX1 inst_cellmath__63_0_I2194 (.CO(N6054), .S(N5867), .A(N6494), .B(N6117), .CI(N5978));
ADDFX1 inst_cellmath__63_0_I2195 (.CO(N6432), .S(N6243), .A(N6008), .B(N6356), .CI(N5867));
ADDFX1 inst_cellmath__63_0_I2196 (.CO(inst_cellmath__63__W1[28]), .S(inst_cellmath__63__W0[27]), .A(N6243), .B(N6388), .CI(N5897));
ADDFX1 inst_cellmath__63_0_I2197 (.CO(N6324), .S(N6135), .A(N6574), .B(N2822), .CI(N5823));
ADDFX1 inst_cellmath__63_0_I2198 (.CO(N5838), .S(N6512), .A(N5766), .B(N5738), .CI(N5796));
ADDFX1 inst_cellmath__63_0_I2199 (.CO(N6212), .S(N6026), .A(N6135), .B(N5790), .CI(N6163));
ADDFX1 inst_cellmath__63_0_I2200 (.CO(N5729), .S(N6403), .A(N6544), .B(N6512), .CI(N6026));
ADDFX1 inst_cellmath__63_0_I2201 (.CO(inst_cellmath__63__W1[29]), .S(inst_cellmath__63__W0[28]), .A(N6403), .B(N6054), .CI(N6432));
ADDFX1 inst_cellmath__63_0_I2202 (.CO(N6480), .S(N6289), .A(N6114), .B(N2887), .CI(N6198));
ADDFX1 inst_cellmath__63_0_I2203 (.CO(N5993), .S(N5805), .A(N6171), .B(N6141), .CI(N6324));
ADDFX1 inst_cellmath__63_0_I2204 (.CO(N6369), .S(N6180), .A(N5838), .B(N6289), .CI(N5805));
ADDFX1 inst_cellmath__63_0_I2205 (.CO(inst_cellmath__63__W1[30]), .S(inst_cellmath__63__W0[29]), .A(N6180), .B(N6212), .CI(N5729));
ADDFX1 inst_cellmath__63_0_I2206 (.CO(N6255), .S(N6068), .A(N6520), .B(N2637), .CI(N6577));
ADDFX1 inst_cellmath__63_0_I2207 (.CO(N5771), .S(N6446), .A(N6480), .B(N6547), .CI(N6068));
ADDFX1 inst_cellmath__63_0_I2208 (.CO(inst_cellmath__63__W1[31]), .S(inst_cellmath__63__W0[30]), .A(N6446), .B(N5993), .CI(N6369));
ADDFX1 inst_cellmath__63_0_I2209 (.CO(N6524), .S(N6335), .A(N6059), .B(N2705), .CI(N6085));
ADDFX1 inst_cellmath__63_0_I2210 (.CO(inst_cellmath__63__W1[32]), .S(inst_cellmath__63__W0[31]), .A(N6335), .B(N6255), .CI(N5771));
ADDFX1 inst_cellmath__63_0_I2211 (.CO(inst_cellmath__63__W1[33]), .S(inst_cellmath__63__W0[32]), .A(N6466), .B(N2776), .CI(N6524));
ADDHX1 inst_cellmath__64_0_I2212 (.CO(N7602), .S(N7477), .A(N477), .B(inst_cellmath__63__W0[15]));
XNOR2X1 inst_cellmath__64_0_I2213 (.Y(N7741), .A(N478), .B(inst_cellmath__63__W0[16]));
OR2XL inst_cellmath__64_0_I2214 (.Y(N7876), .A(N478), .B(inst_cellmath__63__W0[16]));
ADDHX1 inst_cellmath__64_0_I2215 (.CO(N7795), .S(N7663), .A(inst_cellmath__63__W1[16]), .B(inst_cellmath__62__W0[16]));
ADDFX1 inst_cellmath__64_0_I2216 (.CO(N7450), .S(N7929), .A(inst_cellmath__63__W0[17]), .B(N479), .CI(inst_cellmath__63__W1[17]));
ADDHX1 inst_cellmath__64_0_I2217 (.CO(N7720), .S(N7579), .A(inst_cellmath__62__W0[17]), .B(inst_cellmath__62__W1[17]));
ADDFX1 inst_cellmath__64_0_I2218 (.CO(N7979), .S(N7846), .A(inst_cellmath__63__W0[18]), .B(N480), .CI(inst_cellmath__63__W1[18]));
ADDHX1 inst_cellmath__64_0_I2219 (.CO(N7637), .S(N7512), .A(inst_cellmath__62__W0[18]), .B(inst_cellmath__62__W1[18]));
ADDFX1 inst_cellmath__64_0_I2220 (.CO(N7909), .S(N7773), .A(inst_cellmath__63__W0[19]), .B(N481), .CI(inst_cellmath__63__W1[19]));
ADDHX1 inst_cellmath__64_0_I2221 (.CO(N7561), .S(N7427), .A(inst_cellmath__62__W0[19]), .B(inst_cellmath__62__W1[19]));
ADDFX1 inst_cellmath__64_0_I2222 (.CO(N7823), .S(N7698), .A(inst_cellmath__63__W0[20]), .B(N482), .CI(inst_cellmath__63__W1[20]));
ADDHX1 inst_cellmath__64_0_I2223 (.CO(N7489), .S(N7959), .A(inst_cellmath__62__W0[20]), .B(inst_cellmath__62__W1[20]));
ADDFX1 inst_cellmath__64_0_I2224 (.CO(N7753), .S(N7612), .A(inst_cellmath__63__W0[21]), .B(N483), .CI(inst_cellmath__63__W1[21]));
ADDHX1 inst_cellmath__64_0_I2225 (.CO(N7408), .S(N7886), .A(inst_cellmath__62__W0[21]), .B(inst_cellmath__62__W1[21]));
ADDFX1 inst_cellmath__64_0_I2226 (.CO(N7673), .S(N7540), .A(inst_cellmath__63__W0[22]), .B(N484), .CI(inst_cellmath__62__W0[22]));
ADDHX1 inst_cellmath__64_0_I2227 (.CO(N7940), .S(N7804), .A(inst_cellmath__63__W1[22]), .B(inst_cellmath__62__W1[22]));
ADDFX1 inst_cellmath__64_0_I2228 (.CO(N7590), .S(N7461), .A(inst_cellmath__62__W0[23]), .B(N485), .CI(inst_cellmath__62__W1[23]));
ADDHX1 inst_cellmath__64_0_I2229 (.CO(N7859), .S(N7730), .A(inst_cellmath__63__W0[23]), .B(inst_cellmath__63__W1[23]));
ADDFX1 inst_cellmath__64_0_I2230 (.CO(N7523), .S(N7988), .A(inst_cellmath__62__W0[24]), .B(N486), .CI(inst_cellmath__62__W1[24]));
ADDHX1 inst_cellmath__64_0_I2231 (.CO(N7783), .S(N7647), .A(inst_cellmath__63__W0[24]), .B(inst_cellmath__63__W1[24]));
ADDHX1 inst_cellmath__64_0_I2233 (.CO(N7709), .S(N7568), .A(inst_cellmath__63__W0[25]), .B(inst_cellmath__63__W1[25]));
ADDHX1 inst_cellmath__64_0_I2235 (.CO(N7624), .S(N7500), .A(inst_cellmath__63__W0[26]), .B(inst_cellmath__63__W1[26]));
ADDHX1 inst_cellmath__64_0_I2237 (.CO(N7548), .S(N7416), .A(inst_cellmath__63__W0[27]), .B(inst_cellmath__63__W1[27]));
ADDHX1 inst_cellmath__64_0_I2239 (.CO(N7474), .S(N7946), .A(inst_cellmath__63__W0[28]), .B(inst_cellmath__63__W1[28]));
ADDHX1 inst_cellmath__64_0_I2241 (.CO(N7996), .S(N7873), .A(inst_cellmath__63__W0[29]), .B(inst_cellmath__63__W1[29]));
ADDHX1 inst_cellmath__64_0_I2243 (.CO(N7927), .S(N7791), .A(inst_cellmath__63__W0[30]), .B(inst_cellmath__63__W1[30]));
ADDHX1 inst_cellmath__64_0_I2245 (.CO(N7843), .S(N7716), .A(inst_cellmath__63__W0[31]), .B(inst_cellmath__63__W1[31]));
ADDHX1 inst_cellmath__64_0_I2247 (.CO(N7770), .S(N7634), .A(inst_cellmath__63__W0[32]), .B(inst_cellmath__63__W1[32]));
ADDHX1 inst_cellmath__64_0_I2249 (.CO(N7696), .S(N7556), .A(N495), .B(inst_cellmath__63__W1[33]));
NOR4X1 inst_cellmath__64_0_I4936 (.Y(N7895), .A(N6568), .B(N6531), .C(N6299), .D(N6075));
ADDHX1 inst_cellmath__64_0_I2266 (.CO(N7547), .S(N7414), .A(inst_cellmath__63__W1[2]), .B(inst_cellmath__63__W0[2]));
ADDHX1 inst_cellmath__64_0_I2268 (.CO(N7945), .S(N7811), .A(inst_cellmath__63__W1[3]), .B(inst_cellmath__63__W0[3]));
ADDHX1 inst_cellmath__64_0_I2269 (.CO(N7868), .S(N7642), .A(inst_cellmath__63__W0[4]), .B(inst_cellmath__62__W0[4]));
ADDHX1 inst_cellmath__64_0_I2270 (.CO(N7737), .S(N7597), .A(inst_cellmath__63__W1[4]), .B(N7642));
ADDFX1 inst_cellmath__64_0_I2271 (.CO(N7656), .S(N7546), .A(inst_cellmath__62__W1[5]), .B(inst_cellmath__63__W0[5]), .CI(inst_cellmath__62__W0[5]));
ADDFX1 inst_cellmath__64_0_I2272 (.CO(N7528), .S(N7995), .A(N7868), .B(inst_cellmath__63__W1[5]), .CI(N7546));
ADDFX1 inst_cellmath__64_0_I2273 (.CO(N7445), .S(N7444), .A(inst_cellmath__63__W0[6]), .B(inst_cellmath__62__W0[6]), .CI(inst_cellmath__62__W1[6]));
ADDFX1 inst_cellmath__64_0_I2274 (.CO(N7925), .S(N7789), .A(N7656), .B(inst_cellmath__63__W1[6]), .CI(N7444));
ADDFX1 inst_cellmath__64_0_I2275 (.CO(N7839), .S(N7949), .A(inst_cellmath__63__W0[7]), .B(inst_cellmath__62__W0[7]), .CI(inst_cellmath__63__W1[7]));
ADDFX1 inst_cellmath__64_0_I2276 (.CO(N7715), .S(N7574), .A(inst_cellmath__62__W1[7]), .B(N7445), .CI(N7949));
ADDFX1 inst_cellmath__64_0_I2277 (.CO(N7631), .S(N7851), .A(inst_cellmath__62__W0[8]), .B(inst_cellmath__63__W0[8]), .CI(inst_cellmath__63__W1[8]));
ADDFX1 inst_cellmath__64_0_I2278 (.CO(N7506), .S(N7974), .A(N7839), .B(inst_cellmath__62__W1[8]), .CI(N7851));
ADDFX1 inst_cellmath__64_0_I2279 (.CO(N7423), .S(N7757), .A(inst_cellmath__63__W1[9]), .B(inst_cellmath__63__W0[9]), .CI(inst_cellmath__62__W0[9]));
ADDFX1 inst_cellmath__64_0_I2280 (.CO(N7905), .S(N7767), .A(N7631), .B(inst_cellmath__62__W1[9]), .CI(N7757));
ADDFX1 inst_cellmath__64_0_I2281 (.CO(N7819), .S(N7651), .A(inst_cellmath__63__W1[10]), .B(inst_cellmath__63__W0[10]), .CI(inst_cellmath__62__W0[10]));
ADDFX1 inst_cellmath__64_0_I2282 (.CO(N7693), .S(N7555), .A(N7423), .B(inst_cellmath__62__W1[10]), .CI(N7651));
ADDFX1 inst_cellmath__64_0_I2283 (.CO(N7607), .S(N7550), .A(inst_cellmath__63__W1[11]), .B(inst_cellmath__63__W0[11]), .CI(inst_cellmath__62__W0[11]));
ADDFX1 inst_cellmath__64_0_I2284 (.CO(N7481), .S(N7951), .A(N7819), .B(inst_cellmath__62__W1[11]), .CI(N7550));
ADDFX1 inst_cellmath__64_0_I2285 (.CO(N8004), .S(N7452), .A(inst_cellmath__63__W1[12]), .B(inst_cellmath__63__W0[12]), .CI(inst_cellmath__62__W0[12]));
ADDFX1 inst_cellmath__64_0_I2286 (.CO(N7882), .S(N7745), .A(N7452), .B(N7607), .CI(inst_cellmath__62__W1[12]));
ADDFX1 inst_cellmath__64_0_I2287 (.CO(N7800), .S(N7961), .A(inst_cellmath__63__W1[13]), .B(inst_cellmath__63__W0[13]), .CI(inst_cellmath__62__W0[13]));
ADDFX1 inst_cellmath__64_0_I2288 (.CO(N7667), .S(N7534), .A(N8004), .B(inst_cellmath__62__W1[13]), .CI(N7961));
ADDFX1 inst_cellmath__64_0_I2289 (.CO(N7585), .S(N7861), .A(inst_cellmath__63__W1[14]), .B(inst_cellmath__63__W0[14]), .CI(inst_cellmath__62__W0[14]));
ADDFX1 inst_cellmath__64_0_I2290 (.CO(N7456), .S(N7933), .A(N7800), .B(inst_cellmath__62__W1[14]), .CI(N7861));
ADDFX1 inst_cellmath__64_0_I2291 (.CO(N7984), .S(N7762), .A(inst_cellmath__63__W1[15]), .B(N7477), .CI(inst_cellmath__62__W0[15]));
ADDFX1 inst_cellmath__64_0_I2292 (.CO(N7852), .S(N7723), .A(N7585), .B(inst_cellmath__62__W1[15]), .CI(N7762));
ADDFX1 inst_cellmath__64_0_I2293 (.CO(N7778), .S(N7662), .A(N7741), .B(N7602), .CI(inst_cellmath__62__W1[16]));
ADDFX1 inst_cellmath__64_0_I2294 (.CO(N7641), .S(N7515), .A(N7984), .B(N7663), .CI(N7662));
ADDFX1 inst_cellmath__64_0_I2295 (.CO(N7564), .S(N7558), .A(N7929), .B(N7876), .CI(N7795));
ADDFX1 inst_cellmath__64_0_I2296 (.CO(N7431), .S(N7912), .A(N7778), .B(N7579), .CI(N7558));
ADDFX1 inst_cellmath__64_0_I2297 (.CO(N7963), .S(N7459), .A(N7846), .B(N7450), .CI(N7512));
ADDFX1 inst_cellmath__64_0_I2298 (.CO(N7827), .S(N7701), .A(N7564), .B(N7720), .CI(N7459));
ADDFX1 inst_cellmath__64_0_I2299 (.CO(N7758), .S(N7967), .A(N7773), .B(N7979), .CI(N7427));
ADDFX1 inst_cellmath__64_0_I2300 (.CO(N7619), .S(N7492), .A(N7963), .B(N7637), .CI(N7967));
ADDFX1 inst_cellmath__64_0_I2301 (.CO(N7543), .S(N7871), .A(N7698), .B(N7909), .CI(N7561));
ADDFX1 inst_cellmath__64_0_I2302 (.CO(N7412), .S(N7891), .A(N7758), .B(N7959), .CI(N7871));
ADDFX1 inst_cellmath__64_0_I2303 (.CO(N7943), .S(N7769), .A(N7612), .B(N7823), .CI(N7886));
ADDFX1 inst_cellmath__64_0_I2304 (.CO(N7808), .S(N7678), .A(N7543), .B(N7489), .CI(N7769));
ADDFX1 inst_cellmath__64_0_I2305 (.CO(N7734), .S(N7668), .A(N7804), .B(N7753), .CI(N7540));
ADDFX1 inst_cellmath__64_0_I2306 (.CO(N7595), .S(N7465), .A(N7943), .B(N7408), .CI(N7668));
ADDFX1 inst_cellmath__64_0_I2307 (.CO(N7526), .S(N7566), .A(N7461), .B(N7730), .CI(N7940));
ADDFX1 inst_cellmath__64_0_I2308 (.CO(N7992), .S(N7865), .A(N7734), .B(N7673), .CI(N7566));
ADDFX1 inst_cellmath__64_0_I2309 (.CO(N7922), .S(N7468), .A(N7647), .B(N7988), .CI(N7859));
ADDFX1 inst_cellmath__64_0_I2310 (.CO(N7787), .S(N7652), .A(N7526), .B(N7590), .CI(N7468));
ADDFX1 inst_cellmath__64_0_I2311 (.CO(N7713), .S(N7972), .A(N7523), .B(N487), .CI(N7783));
ADDFX1 inst_cellmath__64_0_I2312 (.CO(N7571), .S(N7440), .A(N7922), .B(N7568), .CI(N7972));
ADDHX1 inst_cellmath__64_0_I2313 (.CO(N7503), .S(N7881), .A(N488), .B(N7500));
ADDFX1 inst_cellmath__64_0_I2314 (.CO(N7971), .S(N7835), .A(N7713), .B(N7709), .CI(N7881));
ADDHX1 inst_cellmath__64_0_I2315 (.CO(N7903), .S(N7776), .A(N489), .B(N7416));
ADDFX1 inst_cellmath__64_0_I2316 (.CO(N7764), .S(N7628), .A(N7503), .B(N7624), .CI(N7776));
ADDHX1 inst_cellmath__64_0_I2317 (.CO(N7690), .S(N7676), .A(N490), .B(N7946));
ADDFX1 inst_cellmath__64_0_I2318 (.CO(N7551), .S(N7420), .A(N7903), .B(N7548), .CI(N7676));
ADDHX1 inst_cellmath__64_0_I2319 (.CO(N7479), .S(N7570), .A(N491), .B(N7873));
ADDFX1 inst_cellmath__64_0_I2320 (.CO(N7948), .S(N7817), .A(N7690), .B(N7474), .CI(N7570));
ADDHX1 inst_cellmath__64_0_I2321 (.CO(N7878), .S(N7478), .A(N492), .B(N7791));
ADDFX1 inst_cellmath__64_0_I2322 (.CO(N7742), .S(N7605), .A(N7479), .B(N7996), .CI(N7478));
ADDHX1 inst_cellmath__64_0_I2323 (.CO(N7665), .S(N7980), .A(N493), .B(N7716));
ADDFX1 inst_cellmath__64_0_I2324 (.CO(N7532), .S(N8001), .A(N7878), .B(N7927), .CI(N7980));
ADDHX1 inst_cellmath__64_0_I2325 (.CO(N7453), .S(N7887), .A(N494), .B(N7634));
ADDFX1 inst_cellmath__64_0_I2326 (.CO(N7931), .S(N7798), .A(N7665), .B(N7843), .CI(N7887));
ADDHX1 inst_cellmath__64_0_I2327 (.CO(N7848), .S(N7785), .A(inst_cellmath__63__W0[33]), .B(N7556));
ADDFX1 inst_cellmath__64_0_I2328 (.CO(N7722), .S(N7581), .A(N7453), .B(N7770), .CI(N7785));
ADDHX1 inst_cellmath__64_0_I2329 (.CO(N7639), .S(N7686), .A(1'B1), .B(N496));
ADDFX1 inst_cellmath__64_0_I2330 (.CO(N7514), .S(N7982), .A(N7848), .B(N7696), .CI(N7686));
XNOR2X1 hap1_A_I4941 (.Y(N7775), .A(N497), .B(N7639));
OR2XL hap1_A_I4942 (.Y(N7911), .A(N497), .B(N7639));
INVXL hap1_A_I13852 (.Y(N7484), .A(N498));
OR2XL hap1_A_I4944 (.Y(N7825), .A(1'B0), .B(N498));
INVXL hap1_A_I13853 (.Y(N7987), .A(N499));
OR2XL hap1_A_I4946 (.Y(N7614), .A(1'B0), .B(N499));
ADDHX1 inst_cellmath__64_0_I2336 (.CO(N7491), .S(N7962), .A(N7825), .B(N7987));
XNOR2X1 hap1_A_I4947 (.Y(N7755), .A(N500), .B(N7614));
OR2XL hap1_A_I4948 (.Y(N7889), .A(N500), .B(N7614));
OR2XL inst_cellmath__64_0_I4923 (.Y(N7790), .A(N3894), .B(a_man[22]));
NOR2XL inst_cellmath__64_0_I2346 (.Y(N7990), .A(N7547), .B(N7811));
NAND2XL inst_cellmath__64_0_I2347 (.Y(N7525), .A(N7547), .B(N7811));
AND2XL inst_cellmath__64_0_I2349 (.Y(N7786), .A(N7945), .B(N7597));
NOR2XL inst_cellmath__64_0_I2350 (.Y(N7921), .A(N7737), .B(N7995));
NAND2XL inst_cellmath__64_0_I2351 (.Y(N7436), .A(N7737), .B(N7995));
AND2XL inst_cellmath__64_0_I2353 (.Y(N7711), .A(N7528), .B(N7789));
NOR2XL inst_cellmath__64_0_I2354 (.Y(N7831), .A(N7925), .B(N7574));
NAND2XL inst_cellmath__64_0_I2355 (.Y(N7969), .A(N7925), .B(N7574));
AND2XL inst_cellmath__64_0_I2357 (.Y(N7625), .A(N7715), .B(N7974));
NOR2XL inst_cellmath__64_0_I2358 (.Y(N7763), .A(N7506), .B(N7767));
NAND2XL inst_cellmath__64_0_I2359 (.Y(N7902), .A(N7506), .B(N7767));
AND2XL inst_cellmath__64_0_I2361 (.Y(N7549), .A(N7905), .B(N7555));
NOR2XL inst_cellmath__64_0_I2362 (.Y(N7688), .A(N7693), .B(N7951));
NAND2XL inst_cellmath__64_0_I2363 (.Y(N7814), .A(N7693), .B(N7951));
AND2XL inst_cellmath__64_0_I2365 (.Y(N7476), .A(N7481), .B(N7745));
NOR2XL inst_cellmath__64_0_I2366 (.Y(N7599), .A(N7882), .B(N7534));
NAND2XL inst_cellmath__64_0_I2367 (.Y(N7739), .A(N7882), .B(N7534));
AND2XL inst_cellmath__64_0_I2369 (.Y(N7997), .A(N7667), .B(N7933));
NAND2XL inst_cellmath__64_0_I4937 (.Y(N7636), .A(N7895), .B(N7414));
AOI21XL inst_cellmath__64_0_I2374 (.Y(N7487), .A0(N7525), .A1(N7636), .B0(N7990));
OAI22XL inst_cellmath__64_0_I4925 (.Y(N7857), .A0(N7786), .A1(N7487), .B0(N7945), .B1(N7597));
AOI21XL inst_cellmath__64_0_I2378 (.Y(N7623), .A0(N7436), .A1(N7857), .B0(N7921));
OAI22XL inst_cellmath__64_0_I4926 (.Y(N7926), .A0(N7711), .A1(N7623), .B0(N7528), .B1(N7789));
AOI21XL inst_cellmath__64_0_I2382 (.Y(N7609), .A0(N7969), .A1(N7926), .B0(N7831));
OAI22XL inst_cellmath__64_0_I4927 (.Y(N7828), .A0(N7625), .A1(N7609), .B0(N7715), .B1(N7974));
AOI21XL inst_cellmath__64_0_I2386 (.Y(N7442), .A0(N7902), .A1(N7828), .B0(N7763));
OAI22XL inst_cellmath__64_0_I4928 (.Y(N7583), .A0(N7549), .A1(N7442), .B0(N7905), .B1(N7555));
AOI21XL inst_cellmath__64_0_I2390 (.Y(N7733), .A0(N7814), .A1(N7583), .B0(N7688));
OAI22XL inst_cellmath__64_0_I4929 (.Y(N7796), .A0(N7476), .A1(N7733), .B0(N7481), .B1(N7745));
AOI21XL inst_cellmath__64_0_I2394 (.Y(N7860), .A0(N7739), .A1(N7796), .B0(N7599));
OAI22XL inst_cellmath__64_0_I4930 (.Y(N7694), .A0(N7997), .A1(N7860), .B0(N7667), .B1(N7933));
XOR2XL inst_cellmath__64_0_I2430 (.Y(N8005), .A(N7641), .B(N7912));
XNOR2X1 inst_cellmath__64_0_I2431 (.Y(N7669), .A(N7431), .B(N7701));
XOR2XL inst_cellmath__64_0_I2432 (.Y(N7934), .A(N7827), .B(N7492));
XNOR2X1 inst_cellmath__64_0_I2433 (.Y(N7586), .A(N7619), .B(N7891));
XOR2XL inst_cellmath__64_0_I2434 (.Y(N7853), .A(N7412), .B(N7678));
XNOR2X1 inst_cellmath__64_0_I2435 (.Y(N7517), .A(N7808), .B(N7465));
XOR2XL inst_cellmath__64_0_I2436 (.Y(N7779), .A(N7595), .B(N7865));
XNOR2X1 inst_cellmath__64_0_I2437 (.Y(N7432), .A(N7992), .B(N7652));
XOR2XL inst_cellmath__64_0_I2438 (.Y(N7703), .A(N7440), .B(N7787));
XNOR2X1 inst_cellmath__64_0_I2439 (.Y(N7964), .A(N7571), .B(N7835));
XOR2XL inst_cellmath__64_0_I2440 (.Y(N7620), .A(N7971), .B(N7628));
XNOR2X1 inst_cellmath__64_0_I2441 (.Y(N7893), .A(N7764), .B(N7420));
XOR2XL inst_cellmath__64_0_I2442 (.Y(N7544), .A(N7551), .B(N7817));
XNOR2X1 inst_cellmath__64_0_I2443 (.Y(N7809), .A(N7605), .B(N7948));
XOR2XL inst_cellmath__64_0_I2444 (.Y(N7467), .A(N8001), .B(N7742));
XNOR2X1 inst_cellmath__64_0_I2445 (.Y(N7736), .A(N7798), .B(N7532));
XOR2XL inst_cellmath__64_0_I2446 (.Y(N7993), .A(N7581), .B(N7931));
XNOR2X1 inst_cellmath__64_0_I2447 (.Y(N7654), .A(N7982), .B(N7722));
XOR2XL inst_cellmath__64_0_I2448 (.Y(N7924), .A(N7775), .B(N7514));
XNOR2X1 inst_cellmath__64_0_I2449 (.Y(N7572), .A(N7911), .B(N7484));
XNOR2X1 inst_cellmath__64_0_I2451 (.Y(N7505), .A(N7491), .B(N7755));
XNOR2X1 inst_cellmath__64_0_I2452 (.Y(N7765), .A(N7889), .B(N7790));
INVXL cmpii_A_I13856 (.Y(N22794), .A(N7456));
INVXL cmpii_A_I13857 (.Y(N22796), .A(N7723));
AND2XL cmpii_A_I13858 (.Y(N22792), .A(N22794), .B(N22796));
OAI22XL cmpii_A_I13859 (.Y(N7552), .A0(N22792), .A1(N7694), .B0(N22794), .B1(N22796));
OR2XL cmpoi_A_I4949 (.Y(N11605), .A(N7852), .B(N7515));
AOI22XL cmpoi_A_I4950 (.Y(N8002), .A0(N7552), .A1(N11605), .B0(N7852), .B1(N7515));
AOI2BB2X1 inst_cellmath__64_0_I2455 (.Y(N7850), .A0N(N7641), .A1N(N7912), .B0(N8002), .B1(N8005));
OAI22XL inst_cellmath__64_0_I2456 (.Y(N7617), .A0(N7669), .A1(N7850), .B0(N7431), .B1(N7701));
AOI2BB2X1 inst_cellmath__64_0_I2457 (.Y(N7991), .A0N(N7827), .A1N(N7492), .B0(N7617), .B1(N7934));
OAI22XL inst_cellmath__64_0_I2458 (.Y(N7689), .A0(N7586), .A1(N7991), .B0(N7619), .B1(N7891));
AOI2BB2X1 inst_cellmath__64_0_I2459 (.Y(N7978), .A0N(N7412), .A1N(N7678), .B0(N7689), .B1(N7853));
OAI22XL inst_cellmath__64_0_I2460 (.Y(N7592), .A0(N7517), .A1(N7978), .B0(N7808), .B1(N7465));
AOI2BB2X1 inst_cellmath__64_0_I2461 (.Y(N7812), .A0N(N7595), .A1N(N7865), .B0(N7592), .B1(N7779));
OAI22XL inst_cellmath__64_0_I2462 (.Y(N7954), .A0(N7432), .A1(N7812), .B0(N7992), .B1(N7652));
AOI2BB2X1 inst_cellmath__64_0_I2463 (.Y(N7495), .A0N(N7440), .A1N(N7787), .B0(N7954), .B1(N7703));
OAI22XL inst_cellmath__64_0_I2464 (.Y(N7554), .A0(N7964), .A1(N7495), .B0(N7571), .B1(N7835));
AOI2BB2X1 inst_cellmath__64_0_I2465 (.Y(N7618), .A0N(N7971), .A1N(N7628), .B0(N7554), .B1(N7620));
OAI22XL inst_cellmath__64_0_I2466 (.Y(N7604), .A0(N7893), .A1(N7618), .B0(N7764), .B1(N7420));
AOI2BB2X1 inst_cellmath__64_0_I2467 (.Y(N7593), .A0N(N7551), .A1N(N7817), .B0(N7604), .B1(N7544));
OAI22XL inst_cellmath__64_0_I2468 (.Y(N7510), .A0(N7809), .A1(N7593), .B0(N7605), .B1(N7948));
AOI2BB2X1 inst_cellmath__64_0_I2469 (.Y(N7415), .A0N(N8001), .A1N(N7742), .B0(N7510), .B1(N7467));
OAI22XL inst_cellmath__64_0_I2470 (.Y(N7854), .A0(N7736), .A1(N7415), .B0(N7798), .B1(N7532));
AOI2BB2X1 inst_cellmath__64_0_I2471 (.Y(N7692), .A0N(N7581), .A1N(N7931), .B0(N7854), .B1(N7993));
OAI22XL inst_cellmath__64_0_I2472 (.Y(N7438), .A0(N7654), .A1(N7692), .B0(N7982), .B1(N7722));
AOI2BB2X1 inst_cellmath__64_0_I2473 (.Y(N7806), .A0N(N7775), .A1N(N7514), .B0(N7438), .B1(N7924));
OAI22XL inst_cellmath__64_0_I2474 (.Y(N7486), .A0(N7572), .A1(N7806), .B0(N7911), .B1(N7484));
NOR2BX1 inst_cellmath__64_0_I2475 (.Y(N7768), .AN(N7962), .B(N7486));
OA22X1 inst_cellmath__64_0_I2476 (.Y(N7970), .A0(N7505), .A1(N7768), .B0(N7491), .B1(N7755));
XNOR2X1 inst_cellmath__64_0_I2479 (.Y(inst_cellmath__64[17]), .A(N8002), .B(N8005));
XNOR2X1 inst_cellmath__64_0_I2480 (.Y(inst_cellmath__64[18]), .A(N7850), .B(N7669));
XNOR2X1 inst_cellmath__64_0_I2481 (.Y(inst_cellmath__64[19]), .A(N7617), .B(N7934));
XNOR2X1 inst_cellmath__64_0_I2482 (.Y(inst_cellmath__64[20]), .A(N7991), .B(N7586));
XNOR2X1 inst_cellmath__64_0_I2483 (.Y(inst_cellmath__64[21]), .A(N7689), .B(N7853));
XNOR2X1 inst_cellmath__64_0_I2484 (.Y(inst_cellmath__64[22]), .A(N7978), .B(N7517));
XNOR2X1 inst_cellmath__64_0_I2485 (.Y(inst_cellmath__64[23]), .A(N7592), .B(N7779));
XNOR2X1 inst_cellmath__64_0_I2486 (.Y(inst_cellmath__64[24]), .A(N7812), .B(N7432));
XNOR2X1 inst_cellmath__64_0_I2487 (.Y(inst_cellmath__64[25]), .A(N7954), .B(N7703));
XNOR2X1 inst_cellmath__64_0_I2488 (.Y(inst_cellmath__64[26]), .A(N7495), .B(N7964));
XNOR2X1 inst_cellmath__64_0_I2489 (.Y(inst_cellmath__64[27]), .A(N7554), .B(N7620));
XNOR2X1 inst_cellmath__64_0_I2490 (.Y(inst_cellmath__64[28]), .A(N7618), .B(N7893));
XNOR2X1 inst_cellmath__64_0_I2491 (.Y(inst_cellmath__64[29]), .A(N7604), .B(N7544));
XNOR2X1 inst_cellmath__64_0_I2492 (.Y(inst_cellmath__64[30]), .A(N7593), .B(N7809));
XNOR2X1 inst_cellmath__64_0_I2493 (.Y(inst_cellmath__64[31]), .A(N7510), .B(N7467));
XNOR2X1 inst_cellmath__64_0_I2494 (.Y(inst_cellmath__64[32]), .A(N7415), .B(N7736));
XNOR2X1 inst_cellmath__64_0_I2495 (.Y(inst_cellmath__64[33]), .A(N7854), .B(N7993));
XNOR2X1 inst_cellmath__64_0_I2496 (.Y(inst_cellmath__64[34]), .A(N7692), .B(N7654));
XNOR2X1 inst_cellmath__64_0_I2497 (.Y(inst_cellmath__64[35]), .A(N7438), .B(N7924));
XNOR2X1 inst_cellmath__64_0_I2498 (.Y(inst_cellmath__64[36]), .A(N7806), .B(N7572));
XNOR2X1 inst_cellmath__64_0_I2499 (.Y(inst_cellmath__64[37]), .A(N7486), .B(N7962));
XNOR2X1 inst_cellmath__64_0_I2500 (.Y(inst_cellmath__64[38]), .A(N7768), .B(N7505));
XNOR2X1 inst_cellmath__64_0_I2501 (.Y(inst_cellmath__64[39]), .A(N7970), .B(N7765));
MX2XL inst_cellmath__68_0_I2502 (.Y(x[0]), .A(inst_cellmath__29), .B(inst_cellmath__64[17]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2503 (.Y(x[1]), .A(inst_cellmath__29), .B(inst_cellmath__64[18]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2504 (.Y(x[2]), .A(inst_cellmath__29), .B(inst_cellmath__64[19]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2505 (.Y(x[3]), .A(inst_cellmath__29), .B(inst_cellmath__64[20]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2506 (.Y(x[4]), .A(inst_cellmath__29), .B(inst_cellmath__64[21]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2507 (.Y(x[5]), .A(inst_cellmath__29), .B(inst_cellmath__64[22]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2508 (.Y(x[6]), .A(inst_cellmath__29), .B(inst_cellmath__64[23]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2509 (.Y(x[7]), .A(inst_cellmath__29), .B(inst_cellmath__64[24]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2510 (.Y(x[8]), .A(inst_cellmath__29), .B(inst_cellmath__64[25]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2511 (.Y(x[9]), .A(inst_cellmath__29), .B(inst_cellmath__64[26]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2512 (.Y(x[10]), .A(inst_cellmath__29), .B(inst_cellmath__64[27]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2513 (.Y(x[11]), .A(inst_cellmath__29), .B(inst_cellmath__64[28]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2514 (.Y(x[12]), .A(inst_cellmath__29), .B(inst_cellmath__64[29]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2515 (.Y(x[13]), .A(inst_cellmath__29), .B(inst_cellmath__64[30]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2516 (.Y(x[14]), .A(inst_cellmath__29), .B(inst_cellmath__64[31]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2517 (.Y(x[15]), .A(inst_cellmath__29), .B(inst_cellmath__64[32]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2518 (.Y(x[16]), .A(inst_cellmath__29), .B(inst_cellmath__64[33]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2519 (.Y(x[17]), .A(inst_cellmath__29), .B(inst_cellmath__64[34]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2520 (.Y(x[18]), .A(inst_cellmath__29), .B(inst_cellmath__64[35]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2521 (.Y(x[19]), .A(inst_cellmath__29), .B(inst_cellmath__64[36]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2522 (.Y(x[20]), .A(inst_cellmath__29), .B(inst_cellmath__64[37]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2523 (.Y(x[21]), .A(inst_cellmath__29), .B(inst_cellmath__64[38]), .S0(inst_cellmath__67));
MX2XL inst_cellmath__68_0_I2524 (.Y(x[22]), .A(inst_cellmath__29), .B(inst_cellmath__64[39]), .S0(inst_cellmath__67));
assign inst_cellmath__19[1] = 1'B1;
assign inst_cellmath__19[2] = 1'B1;
assign inst_cellmath__19[3] = 1'B1;
assign inst_cellmath__19[4] = 1'B1;
assign inst_cellmath__19[5] = 1'B1;
assign inst_cellmath__19[6] = 1'B1;
assign inst_cellmath__19[7] = 1'B1;
assign inst_cellmath__19[8] = 1'B1;
assign inst_cellmath__20[2] = 1'B0;
assign inst_cellmath__20[4] = 1'B0;
assign inst_cellmath__20[6] = 1'B0;
assign inst_cellmath__22[8] = 1'B0;
assign inst_cellmath__51[18] = 1'B1;
assign inst_cellmath__62__W0[0] = 1'B0;
assign inst_cellmath__62__W0[1] = 1'B0;
assign inst_cellmath__62__W0[2] = 1'B0;
assign inst_cellmath__62__W0[3] = 1'B0;
assign inst_cellmath__62__W0[25] = 1'B0;
assign inst_cellmath__62__W0[26] = 1'B0;
assign inst_cellmath__62__W0[27] = 1'B0;
assign inst_cellmath__62__W0[28] = 1'B0;
assign inst_cellmath__62__W0[29] = 1'B0;
assign inst_cellmath__62__W0[30] = 1'B0;
assign inst_cellmath__62__W0[31] = 1'B0;
assign inst_cellmath__62__W0[32] = 1'B0;
assign inst_cellmath__62__W0[33] = 1'B0;
assign inst_cellmath__62__W0[34] = 1'B0;
assign inst_cellmath__62__W0[35] = 1'B0;
assign inst_cellmath__62__W0[36] = 1'B0;
assign inst_cellmath__62__W0[37] = 1'B0;
assign inst_cellmath__62__W0[38] = 1'B0;
assign inst_cellmath__62__W0[39] = 1'B0;
assign inst_cellmath__62__W1[0] = 1'B0;
assign inst_cellmath__62__W1[1] = 1'B0;
assign inst_cellmath__62__W1[2] = 1'B0;
assign inst_cellmath__62__W1[3] = 1'B0;
assign inst_cellmath__62__W1[4] = 1'B0;
assign inst_cellmath__62__W1[25] = 1'B0;
assign inst_cellmath__62__W1[26] = 1'B0;
assign inst_cellmath__62__W1[27] = 1'B0;
assign inst_cellmath__62__W1[28] = 1'B0;
assign inst_cellmath__62__W1[29] = 1'B0;
assign inst_cellmath__62__W1[30] = 1'B0;
assign inst_cellmath__62__W1[31] = 1'B0;
assign inst_cellmath__62__W1[32] = 1'B0;
assign inst_cellmath__62__W1[33] = 1'B0;
assign inst_cellmath__62__W1[34] = 1'B0;
assign inst_cellmath__62__W1[35] = 1'B0;
assign inst_cellmath__62__W1[36] = 1'B0;
assign inst_cellmath__62__W1[37] = 1'B0;
assign inst_cellmath__62__W1[38] = 1'B0;
assign inst_cellmath__62__W1[39] = 1'B0;
assign inst_cellmath__63__W0[0] = 1'B0;
assign inst_cellmath__63__W0[1] = 1'B0;
assign inst_cellmath__63__W0[34] = 1'B1;
assign inst_cellmath__63__W0[35] = 1'B1;
assign inst_cellmath__63__W0[36] = 1'B1;
assign inst_cellmath__63__W0[37] = 1'B1;
assign inst_cellmath__63__W0[38] = 1'B1;
assign inst_cellmath__63__W0[39] = 1'B1;
assign inst_cellmath__63__W1[0] = 1'B0;
assign inst_cellmath__63__W1[1] = 1'B0;
assign inst_cellmath__63__W1[34] = 1'B0;
assign inst_cellmath__63__W1[35] = 1'B0;
assign inst_cellmath__63__W1[36] = 1'B0;
assign inst_cellmath__63__W1[37] = 1'B0;
assign inst_cellmath__63__W1[38] = 1'B0;
assign inst_cellmath__63__W1[39] = 1'B0;
assign inst_cellmath__64[0] = 1'B0;
assign inst_cellmath__64[1] = 1'B0;
assign inst_cellmath__64[2] = 1'B0;
assign inst_cellmath__64[3] = 1'B0;
assign inst_cellmath__64[4] = 1'B0;
assign inst_cellmath__64[5] = 1'B0;
assign inst_cellmath__64[6] = 1'B0;
assign inst_cellmath__64[7] = 1'B0;
assign inst_cellmath__64[8] = 1'B0;
assign inst_cellmath__64[9] = 1'B0;
assign inst_cellmath__64[10] = 1'B0;
assign inst_cellmath__64[11] = 1'B0;
assign inst_cellmath__64[12] = 1'B0;
assign inst_cellmath__64[13] = 1'B0;
assign inst_cellmath__64[14] = 1'B0;
assign inst_cellmath__64[15] = 1'B0;
assign inst_cellmath__64[16] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  ubT5QgjWrhA= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



