/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:06:59 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51;
wire [24:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2600,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2617,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2641,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2717,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2828,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795;
wire N11500,N11504,N11506,N11667,N11672,N11677,N11682 
	,N11687,N11692,N11697,N11702,N11707,N11712,N11717,N11722 
	,N11788,N11798,N11806,N11814,N11822,N11830,N11838,N11846 
	,N11854,N11862,N11886,N11937,N11941,N11966,N12003,N12007 
	,N12042,N12044,N12077,N12085,N12087,N12089,N12122,N12130 
	,N12132,N12167,N12169,N12175,N12177,N12183,N12218,N12220 
	,N12238,N12240,N12242,N12277,N12279,N12285,N12289,N12293 
	,N12295,N12297,N12325,N12327,N12363,N12365,N12383,N12413 
	,N12415,N12421,N12423,N12429,N12435,N12443,N12445,N12447 
	,N12480,N12482,N12488,N12490,N12492,N12496,N12498,N12500 
	,N12504,N12506,N12508,N12512,N12514,N12516,N12529,N12542 
	,N12544,N12550,N12552,N12554,N12560,N12562,N12564,N12567 
	,N12578,N12580,N12582,N12585,N12587,N12589,N12591,N12605 
	,N12607,N12609,N12613,N12618,N12625,N12627,N13149,N13150 
	,N13151,N13152,N13153,N13154,N13155,N13156,N13164,N13166 
	,N13167,N13170,N13172,N13174,N13178,N13180,N13181,N13182 
	,N13202,N13204,N13205,N13209,N13212,N13215,N13229,N13232 
	,N13234,N13236,N13238,N13241,N13242,N13246,N13248,N13250 
	,N13251,N13254,N13256,N13259,N13263,N13264,N13266,N13267 
	,N13268,N13269,N13271,N13273,N13274,N13277,N13279,N13281 
	,N13318,N13319,N13322,N13326,N13329,N13330,N13337,N13353 
	,N13354,N13356,N13358,N13359,N13360,N13362,N13364,N13366 
	,N13368,N13370,N13371,N13373,N13376,N13378,N13380,N13382 
	,N13385,N13389,N13391,N13392,N13395,N13400,N13436,N13440 
	,N13443,N13445,N13447,N13450,N13452,N13455,N13457,N13459 
	,N13460,N13461,N13463,N13464,N13466,N13468,N13470,N13472 
	,N13474,N13476,N13478,N13479,N13482,N13484,N13486,N13518 
	,N13521,N13530,N13542,N13543,N13546,N13548,N13550,N13551 
	,N13553,N13556,N13557,N13562,N13564,N13566,N13568,N13570 
	,N13571,N13573,N13575,N13577,N13579,N13581,N13583,N13586 
	,N13588,N13590,N13591,N13626,N13628,N13630,N13632,N13634 
	,N13636,N13639,N13642,N13645,N13647,N13649,N13650,N13651 
	,N13653,N13655,N13659,N13661,N13663,N13665,N13667,N13668 
	,N13671;
reg x_reg_22__retimed_I7284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7284_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14];
	end
assign N12627 = x_reg_22__retimed_I7284_QOUT;
reg x_reg_22__retimed_I7283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7283_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13];
	end
assign N12625 = x_reg_22__retimed_I7283_QOUT;
reg x_reg_22__retimed_I7278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7278_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648;
	end
assign N12609 = x_reg_22__retimed_I7278_QOUT;
reg x_reg_22__retimed_I7277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7277_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832;
	end
assign N12607 = x_reg_22__retimed_I7277_QOUT;
reg x_reg_22__retimed_I7276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7276_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11];
	end
assign N12605 = x_reg_22__retimed_I7276_QOUT;
reg x_reg_22__retimed_I7272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7272_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564;
	end
assign N12591 = x_reg_22__retimed_I7272_QOUT;
reg x_reg_22__retimed_I7271_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7271_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570;
	end
assign N12589 = x_reg_22__retimed_I7271_QOUT;
reg x_reg_22__retimed_I7270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7270_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919;
	end
assign N12587 = x_reg_22__retimed_I7270_QOUT;
reg x_reg_22__retimed_I7269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7269_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800;
	end
assign N12585 = x_reg_22__retimed_I7269_QOUT;
reg x_reg_22__retimed_I7268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7268_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13];
	end
assign N12582 = x_reg_22__retimed_I7268_QOUT;
reg x_reg_22__retimed_I7267_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7267_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13];
	end
assign N12580 = x_reg_22__retimed_I7267_QOUT;
reg x_reg_22__retimed_I7266_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7266_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13];
	end
assign N12578 = x_reg_22__retimed_I7266_QOUT;
reg x_reg_22__retimed_I7262_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7262_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703;
	end
assign N12567 = x_reg_22__retimed_I7262_QOUT;
reg x_reg_22__retimed_I7261_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7261_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12];
	end
assign N12564 = x_reg_22__retimed_I7261_QOUT;
reg x_reg_22__retimed_I7260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7260_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550;
	end
assign N12562 = x_reg_22__retimed_I7260_QOUT;
reg x_reg_22__retimed_I7259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7259_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622;
	end
assign N12560 = x_reg_22__retimed_I7259_QOUT;
reg x_reg_22__retimed_I7258_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7258_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359;
	end
assign N12554 = x_reg_22__retimed_I7258_QOUT;
reg x_reg_22__retimed_I7257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7257_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265;
	end
assign N12552 = x_reg_22__retimed_I7257_QOUT;
reg x_reg_22__retimed_I7256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7256_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209;
	end
assign N12550 = x_reg_22__retimed_I7256_QOUT;
reg x_reg_22__retimed_I7254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7254_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14];
	end
assign N12544 = x_reg_22__retimed_I7254_QOUT;
reg x_reg_22__retimed_I7253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7253_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14];
	end
assign N12542 = x_reg_22__retimed_I7253_QOUT;
reg x_reg_22__retimed_I7248_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7248_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024;
	end
assign N12529 = x_reg_22__retimed_I7248_QOUT;
reg x_reg_22__retimed_I7244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7244_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295;
	end
assign N12516 = x_reg_22__retimed_I7244_QOUT;
reg x_reg_22__retimed_I7243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7243_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283;
	end
assign N12514 = x_reg_22__retimed_I7243_QOUT;
reg x_reg_22__retimed_I7242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7242_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149;
	end
assign N12512 = x_reg_22__retimed_I7242_QOUT;
reg x_reg_22__retimed_I7241_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7241_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275;
	end
assign N12508 = x_reg_22__retimed_I7241_QOUT;
reg x_reg_22__retimed_I7240_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7240_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075;
	end
assign N12506 = x_reg_22__retimed_I7240_QOUT;
reg x_reg_22__retimed_I7239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7239_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128;
	end
assign N12504 = x_reg_22__retimed_I7239_QOUT;
reg x_reg_22__retimed_I7238_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7238_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351;
	end
assign N12500 = x_reg_22__retimed_I7238_QOUT;
reg x_reg_22__retimed_I7237_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7237_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257;
	end
assign N12498 = x_reg_22__retimed_I7237_QOUT;
reg x_reg_22__retimed_I7236_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7236_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203;
	end
assign N12496 = x_reg_22__retimed_I7236_QOUT;
reg x_reg_22__retimed_I7235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7235_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184;
	end
assign N12492 = x_reg_22__retimed_I7235_QOUT;
reg x_reg_22__retimed_I7234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7234_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378;
	end
assign N12490 = x_reg_22__retimed_I7234_QOUT;
reg x_reg_22__retimed_I7233_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7233_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092;
	end
assign N12488 = x_reg_22__retimed_I7233_QOUT;
reg x_reg_22__retimed_I7231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7231_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15];
	end
assign N12482 = x_reg_22__retimed_I7231_QOUT;
reg x_reg_22__retimed_I7230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7230_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487;
	end
assign N12480 = x_reg_22__retimed_I7230_QOUT;
reg x_reg_22__retimed_I7218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7218_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167;
	end
assign N12447 = x_reg_22__retimed_I7218_QOUT;
reg x_reg_22__retimed_I7217_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7217_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358;
	end
assign N12445 = x_reg_22__retimed_I7217_QOUT;
reg x_reg_22__retimed_I7216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7216_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343;
	end
assign N12443 = x_reg_22__retimed_I7216_QOUT;
reg x_reg_22__retimed_I7213_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7213_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090;
	end
assign N12435 = x_reg_22__retimed_I7213_QOUT;
reg x_reg_22__retimed_I7211_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7211_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16];
	end
assign N12429 = x_reg_22__retimed_I7211_QOUT;
reg x_reg_22__retimed_I7209_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7209_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083;
	end
assign N12423 = x_reg_22__retimed_I7209_QOUT;
reg x_reg_22__retimed_I7208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7208_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223;
	end
assign N12421 = x_reg_22__retimed_I7208_QOUT;
reg x_reg_22__retimed_I7206_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7206_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757;
	end
assign N12415 = x_reg_22__retimed_I7206_QOUT;
reg x_reg_22__retimed_I7205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7205_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618;
	end
assign N12413 = x_reg_22__retimed_I7205_QOUT;
reg x_reg_22__retimed_I7194_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7194_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155;
	end
assign N12383 = x_reg_22__retimed_I7194_QOUT;
reg x_reg_22__retimed_I7188_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7188_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945;
	end
assign N12365 = x_reg_22__retimed_I7188_QOUT;
reg x_reg_22__retimed_I7187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7187_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890;
	end
assign N12363 = x_reg_22__retimed_I7187_QOUT;
reg x_reg_22__retimed_I7174_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7174_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864;
	end
assign N12327 = x_reg_22__retimed_I7174_QOUT;
reg x_reg_22__retimed_I7173_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7173_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457;
	end
assign N12325 = x_reg_22__retimed_I7173_QOUT;
reg x_reg_22__retimed_I7163_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7163_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288;
	end
assign N12297 = x_reg_22__retimed_I7163_QOUT;
reg x_reg_22__retimed_I7162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7162_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317;
	end
assign N12295 = x_reg_22__retimed_I7162_QOUT;
reg x_reg_22__retimed_I7161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7161_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143;
	end
assign N12293 = x_reg_22__retimed_I7161_QOUT;
reg x_reg_22__retimed_I7160_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7160_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213;
	end
assign N12289 = x_reg_22__retimed_I7160_QOUT;
reg x_reg_22__retimed_I7158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7158_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228;
	end
assign N12285 = x_reg_22__retimed_I7158_QOUT;
reg x_reg_22__retimed_I7156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7156_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787;
	end
assign N12279 = x_reg_22__retimed_I7156_QOUT;
reg x_reg_22__retimed_I7155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7155_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001;
	end
assign N12277 = x_reg_22__retimed_I7155_QOUT;
reg x_reg_22__retimed_I7143_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7143_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392;
	end
assign N12242 = x_reg_22__retimed_I7143_QOUT;
reg x_reg_22__retimed_I7142_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7142_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272;
	end
assign N12240 = x_reg_22__retimed_I7142_QOUT;
reg x_reg_22__retimed_I7141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7141_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244;
	end
assign N12238 = x_reg_22__retimed_I7141_QOUT;
reg x_reg_22__retimed_I7135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7135_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709;
	end
assign N12220 = x_reg_22__retimed_I7135_QOUT;
reg x_reg_22__retimed_I7134_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7134_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924;
	end
assign N12218 = x_reg_22__retimed_I7134_QOUT;
reg x_reg_22__retimed_I7122_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7122_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22];
	end
assign N12183 = x_reg_22__retimed_I7122_QOUT;
reg x_reg_22__retimed_I7120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7120_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22];
	end
assign N12177 = x_reg_22__retimed_I7120_QOUT;
reg x_reg_22__retimed_I7119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7119_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484;
	end
assign N12175 = x_reg_22__retimed_I7119_QOUT;
reg x_reg_22__retimed_I7117_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7117_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627;
	end
assign N12169 = x_reg_22__retimed_I7117_QOUT;
reg x_reg_22__retimed_I7116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7116_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838;
	end
assign N12167 = x_reg_22__retimed_I7116_QOUT;
reg x_reg_22__retimed_I7104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7104_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23];
	end
assign N12132 = x_reg_22__retimed_I7104_QOUT;
reg x_reg_22__retimed_I7103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7103_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485;
	end
assign N12130 = x_reg_22__retimed_I7103_QOUT;
reg x_reg_22__retimed_I7100_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7100_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767;
	end
assign N12122 = x_reg_22__retimed_I7100_QOUT;
reg x_reg_22__retimed_I7089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7089_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24];
	end
assign N12089 = x_reg_22__retimed_I7089_QOUT;
reg x_reg_22__retimed_I7088_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7088_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24];
	end
assign N12087 = x_reg_22__retimed_I7088_QOUT;
reg x_reg_22__retimed_I7087_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7087_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486;
	end
assign N12085 = x_reg_22__retimed_I7087_QOUT;
reg x_reg_22__retimed_I7084_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7084_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741;
	end
assign N12077 = x_reg_22__retimed_I7084_QOUT;
reg x_reg_22__retimed_I7073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7073_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874;
	end
assign N12044 = x_reg_22__retimed_I7073_QOUT;
reg x_reg_22__retimed_I7072_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7072_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659;
	end
assign N12042 = x_reg_22__retimed_I7072_QOUT;
reg x_reg_22__retimed_I7060_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7060_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795;
	end
assign N12007 = x_reg_22__retimed_I7060_QOUT;
reg x_reg_22__retimed_I7058_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7058_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487;
	end
assign N12003 = x_reg_22__retimed_I7058_QOUT;
reg x_reg_22__retimed_I7045_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7045_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585;
	end
assign N11966 = x_reg_22__retimed_I7045_QOUT;
reg x_reg_22__retimed_I7037_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7037_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982;
	end
assign N11941 = x_reg_22__retimed_I7037_QOUT;
reg x_reg_22__retimed_I7035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7035_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719;
	end
assign N11937 = x_reg_22__retimed_I7035_QOUT;
reg x_reg_22__retimed_I7017_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7017_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638;
	end
assign N11886 = x_reg_22__retimed_I7017_QOUT;
reg x_reg_22__retimed_I7008_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7008_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976;
	end
assign N11862 = x_reg_22__retimed_I7008_QOUT;
reg x_reg_22__retimed_I7005_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7005_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683;
	end
assign N11854 = x_reg_22__retimed_I7005_QOUT;
reg x_reg_22__retimed_I7002_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7002_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009;
	end
assign N11846 = x_reg_22__retimed_I7002_QOUT;
reg x_reg_22__retimed_I6999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6999_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716;
	end
assign N11838 = x_reg_22__retimed_I6999_QOUT;
reg x_reg_22__retimed_I6996_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6996_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418;
	end
assign N11830 = x_reg_22__retimed_I6996_QOUT;
reg x_reg_22__retimed_I6993_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6993_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749;
	end
assign N11822 = x_reg_22__retimed_I6993_QOUT;
reg x_reg_22__retimed_I6990_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6990_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452;
	end
assign N11814 = x_reg_22__retimed_I6990_QOUT;
reg x_reg_22__retimed_I6987_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6987_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781;
	end
assign N11806 = x_reg_22__retimed_I6987_QOUT;
reg x_reg_22__retimed_I6984_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6984_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492;
	end
assign N11798 = x_reg_22__retimed_I6984_QOUT;
reg x_reg_22__retimed_I6981_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6981_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985;
	end
assign N11788 = x_reg_22__retimed_I6981_QOUT;
reg x_reg_11__retimed_I6955_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6955_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896;
	end
assign N11722 = x_reg_11__retimed_I6955_QOUT;
reg x_reg_12__retimed_I6953_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I6953_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546;
	end
assign N11717 = x_reg_12__retimed_I6953_QOUT;
reg x_reg_13__retimed_I6951_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I6951_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813;
	end
assign N11712 = x_reg_13__retimed_I6951_QOUT;
reg x_reg_14__retimed_I6949_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6949_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465;
	end
assign N11707 = x_reg_14__retimed_I6949_QOUT;
reg x_reg_15__retimed_I6947_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I6947_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735;
	end
assign N11702 = x_reg_15__retimed_I6947_QOUT;
reg x_reg_16__retimed_I6945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I6945_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006;
	end
assign N11697 = x_reg_16__retimed_I6945_QOUT;
reg x_reg_17__retimed_I6943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6943_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654;
	end
assign N11692 = x_reg_17__retimed_I6943_QOUT;
reg x_reg_18__retimed_I6941_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I6941_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929;
	end
assign N11687 = x_reg_18__retimed_I6941_QOUT;
reg x_reg_19__retimed_I6939_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6939_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580;
	end
assign N11682 = x_reg_19__retimed_I6939_QOUT;
reg x_reg_20__retimed_I6937_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6937_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983;
	end
assign N11677 = x_reg_20__retimed_I6937_QOUT;
reg x_reg_21__retimed_I6935_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6935_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503;
	end
assign N11672 = x_reg_21__retimed_I6935_QOUT;
reg x_reg_22__retimed_I6933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6933_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772;
	end
assign N11667 = x_reg_22__retimed_I6933_QOUT;
reg x_reg_22__retimed_I6864_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6864_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29;
	end
assign N11506 = x_reg_22__retimed_I6864_QOUT;
assign N13149 = !N11506;
assign N13150 = !N13149;
reg x_reg_22__retimed_I6863_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6863_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67;
	end
assign N11504 = x_reg_22__retimed_I6863_QOUT;
assign N13151 = !N11504;
assign N13156 = !N13151;
assign N13155 = !N13151;
assign N13154 = !N13151;
assign N13153 = !N13151;
reg x_reg_22__retimed_I6861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6861_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795;
	end
assign N11500 = x_reg_22__retimed_I6861_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353 = !(a_exp[7] & a_exp[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355 = ((a_exp[4] & a_exp[3]) & a_exp[2]) & a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743 = !((a_exp[6] & a_exp[5]) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393 = !(((a_man[0] | a_man[1]) | a_man[2]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 = !(a_man[18] | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402 = !((((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381) | a_man[16]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408) | a_man[15]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0] | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1] = !a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0] = !a_exp[0];
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2] = (!a_exp[2]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3] = !a_exp[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457 = !(a_exp[2] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5] = !a_exp[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451 = !(a_exp[4] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6] = (!a_exp[6]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7] = !a_exp[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444 = !(a_exp[6] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4] = (!a_exp[4]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483 = !((((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448 = ((float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427 = !a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 = !a_man[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 = !a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 = !a_man[20];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 = !a_man[18];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 = !(a_man[16] & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 = !a_man[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 = !a_man[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 = !(a_man[17] & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 = !(a_man[17] | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (a_man[19] & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054 = !(a_man[19] | a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[16]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 = !(a_man[17] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 = !((a_man[17] & a_man[16]) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783} = {1'B0, 1'B1} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] = !a_man[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589 & a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 = !a_man[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 = !a_man[13];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16] = !(a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[18] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637 = !a_man[12];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848 | a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888 = !a_man[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 = !a_man[10];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747 = !a_man[9];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648 = !a_man[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 = !a_man[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[18] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 = !a_man[6];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698 = !a_man[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631 = !a_man[4];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 = !a_man[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 = !a_man[2];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 = !a_man[0];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 = !a_man[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 = a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2801 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2821 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2600 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2821} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2801} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2600};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign N13667 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719;
assign N13630 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign {N13649, N13639} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663, N13661} = {1'B0, N13630} + {1'B0, N13667} + {1'B0, N13649};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2649, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2581} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2792, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2717} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2686, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2617} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2581} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2686} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2717};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2617};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614, N13556} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790;
assign {N13590, N13579} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754, N13550} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724} + {1'B0, N13590};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2677, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2608} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647};
assign {N13583, N13570} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2677} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896, N13542} = {1'B0, N13556} + {1'B0, N13583} + {1'B0, N13550};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702, N13440} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2760, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2688} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign {N13474, N13459} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846, N13486} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856} + {1'B0, N13474} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2688};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595};
assign {N13466, N13452} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660, N13478} = {1'B0, N13466} + {1'B0, N13440} + {1'B0, N13486};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11756 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626};
assign {N13445, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586) | (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800);
assign {N13457, N13447} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721};
assign {N13484, N13472} = {1'B0, N13459} + {1'B0, N13457} + {1'B0, N13452};
assign N13443 = !N13484;
assign N13468 = !N13443;
assign N13479 = !((N13478 & N13443) | ((!N13478) & N13468));
assign {N13464, N13450} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615} + {1'B0, N13447};
assign N13476 = N13464 ^ N13472;
assign N13455 = N13445 & N13450;
assign N13470 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797);
assign N13482 = ((!N13445) & (!N13450)) | ((!N13455) & (!N13470));
assign N13461 = !N13472;
assign N13436 = !N13464;
assign N13463 = !((N13436 & N13461) | (N13476 & N13482));
assign N13460 = N13484 | N13478;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576 = ((!N13479) & (!N13463)) | (!N13460);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11758 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576);
assign {N13577, N13564} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794};
assign {N13548, N13588} = {1'B0, N13577} + {1'B0, N13579} + {1'B0, N13570};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795 = N13548 ^ N13542;
assign {N13581, N13568} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2760} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2608} + {1'B0, N13564};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652 = N13581 ^ N13588;
assign N13553 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583 ^ N13568;
assign N13562 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11756 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11758);
assign N13575 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583 | N13568);
assign N13557 = !((N13562 & N13553) | N13575);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871 = (N13562 & N13553) | N13575;
assign N13571 = !N13588;
assign N13543 = !N13581;
assign N13546 = !(N13581 | N13588);
assign N13586 = !(N13557 | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652));
assign N13573 = !(N13546 | N13586);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749 = (N13543 & N13571) | N13586;
assign N13566 = !(N13548 | N13542);
assign N13551 = !(N13573 | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795));
assign N13591 = !(N13566 | N13551);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766 = !N13591;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2828 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2828;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2641 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858);
assign {N13642, N13634} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711};
assign N13655 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708;
assign {N13628, N13665} = {1'B0, N13655} + {1'B0, N13642} + {1'B0, N13639};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813 = N13661 ^ N13628;
assign {N13659, N13647} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2649} + {1'B0, N13634} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2792};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667 = N13659 ^ N13665;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852 = N13647 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2641;
assign N13653 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606 | N13647);
assign N13636 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852) | N13653);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852) | N13653;
assign N13650 = !N13665;
assign N13671 = !N13659;
assign N13626 = !(N13665 | N13659);
assign N13663 = !(N13636 | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667));
assign N13651 = !(N13626 | N13663);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601 = (N13671 & N13650) | N13663;
assign N13645 = !(N13661 | N13628);
assign N13632 = !(N13651 | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813));
assign N13668 = !(N13645 | N13632);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634 = !N13668;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2881 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2881;
assign N13530 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809);
assign N13518 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769) | N13530;
assign N13521 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176 = N13521 ^ N13518;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23] = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917 = !(a_man[21] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010} = {1'B0, N12085} + {1'B0, N12087} + {1'B0, N12089};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332 = !(a_man[16] & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722, N13370} = {1'B0, N12003} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530} + {1'B0, N12007};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853} = {1'B0, N11937} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722} + {1'B0, N11941};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]};
assign {N13400, N13391} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010} + {1'B0, N12042} + {1'B0, N12044};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589, N13364} = {1'B0, N11966} + {1'B0, N13400} + {1'B0, N13370};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]} = {1'B0, N12238} + {1'B0, N12240} + {1'B0, N12242};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552} = {1'B0, N12175} + {1'B0, N12177} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]} = {1'B0, N12293} + {1'B0, N12295} + {1'B0, N12297};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817} = {1'B0, N12183} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770} = {1'B0, N12122} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299} = {1'B0, N12443} + {1'B0, N12445} + {1'B0, N12447};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]} = {1'B0, N12285} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376} + {1'B0, N12289};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868} = {1'B0, N12167} + {1'B0, N12169} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370} = {1'B0, N12504} + {1'B0, N12506} + {1'B0, N12508};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239} = {1'B0, N12516} + {1'B0, N12512} + {1'B0, N12514};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]} = {1'B0, N12435} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]} = {1'B0, N12383} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557, N13256} = {1'B0, N12218} + {1'B0, N12220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497, N13281} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]};
assign {N13259, N13248} = {1'B0, N12277} + {1'B0, N12279} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415, N13273} = {1'B0, N13281} + {1'B0, N13259} + {1'B0, N13256};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]} = {1'B0, N12421} + {1'B0, N12423} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]} = {1'B0, N12488} + {1'B0, N12490} + {1'B0, N12492};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675} = {1'B0, N12429} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655} = {1'B0, N12363} + {1'B0, N12365} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]} = {1'B0, N12496} + {1'B0, N12498} + {1'B0, N12500};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763} = {1'B0, N12413} + {1'B0, N12415} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]} = {1'B0, N12550} + {1'B0, N12552} + {1'B0, N12554};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861} = {1'B0, N12480} + {1'B0, N12482} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964} = {1'B0, N12542} + {1'B0, N12544} + {1'B0, N12627};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442} = {1'B0, N12578} + {1'B0, N12580} + {1'B0, N12582};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545} = {1'B0, N12625} + {1'B0, N12529} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971} = {1'B0, N12605} + {1'B0, N12607} + {1'B0, N12609};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761} = {1'B0, N12560} + {1'B0, N12562} + {1'B0, N12564};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826 = !(N12567 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948 = ((!N12591) & (!N12585)) | ((!N12587) & (!N12589));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699 = !(N12567 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615;
assign N12613 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419) | (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558 = !N12613;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733) & (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524) & (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927;
assign {N13254, N13241} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]};
assign {N13279, N13263} = {1'B0, N12325} + {1'B0, N12327} + {1'B0, N13241};
assign {N13246, N13236} = {1'B0, N13279} + {1'B0, N13254} + {1'B0, N13248};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593 = N13246 ^ N13273;
assign {N13229, N13271} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730} + {1'B0, N13263};
assign N13274 = !N13229;
assign N13251 = !(N13274 | N13236);
assign N13232 = !N13251;
assign N13266 = !N13229;
assign N13238 = !(N13266 & N13236);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940 = N13236 ^ N13229;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439 ^ N13271;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590);
assign N13277 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439 | N13271;
assign N13234 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462 = (!N13277) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668);
assign N13242 = !N13236;
assign N13264 = !(N13229 | N13236);
assign N13269 = !((N13232 & N13238) | (N13277 & N13234));
assign N13250 = !N13269;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500 = (!N13250) | (N13242 & N13274);
assign N13268 = N13246 | N13273;
assign N13267 = ((!N13269) & (!N13264)) | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798 = !(N13268 & N13267);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821;
assign {N13395, N13385} = {1'B0, N12130} + {1'B0, N12132} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23]};
assign {N13368, N13353} = {1'B0, N12077} + {1'B0, N13385} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686};
assign {N13389, N13380} = {1'B0, N13395} + {1'B0, N13368} + {1'B0, N13391};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704 = N13364 ^ N13389;
assign {N13373, N13362} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744} + {1'B0, N13353};
assign N13371 = !N13380;
assign N13376 = !(N13373 & N13371);
assign N13356 = !N13373;
assign N13382 = !(N13380 & N13356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430 = N13373 ^ N13380;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782 = N13362 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756);
assign N13366 = N13362 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610;
assign N13378 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847 = (!N13366) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979);
assign N13354 = !(N13373 | N13380);
assign N13360 = !((N13376 & N13382) | (N13366 & N13378));
assign N13392 = !N13360;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996 = (!N13392) | (N13371 & N13356);
assign N13359 = N13364 | N13389;
assign N13358 = ((!N13360) & (!N13354)) | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794 = !(N13359 & N13358);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623 = N11886 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794);
assign N13337 = N11886 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992;
assign N13329 = !N13337;
assign N13319 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623) | N13329);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579 = (!N13337) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856);
assign N13318 = !N11722;
assign N13326 = !(N13318 | N13319);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567 = (!N11862) | (N11722 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579);
assign N13322 = !N11862;
assign N13330 = ((!N13326) & (!N13322)) | (!N11717);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820 = !(N11854 & N13330);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728 = (!N11846) | (N11712 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911 = (!N11838) | (N11707 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736 = (!N11830) | (N11702 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831 = (!N11822) | (N11697 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736);
assign N13204 = !N11814;
assign N13205 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831 & N11692) | N13204);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588 = (!N11814) | (N11692 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831);
assign N13209 = !N11687;
assign N13212 = !(N13209 | N13205);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608 = (!N11806) | (N11687 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588);
assign N13202 = !N11806;
assign N13215 = ((!N13212) & (!N13202)) | (!N11682);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899 = !(N11798 & N13215);
assign N12618 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899 | (!N11677));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499);
assign N13167 = !N11788;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834 = !N12618;
assign N13180 = !(N11672 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834);
assign N13172 = !N11667;
assign N13181 = !((N13180 & N13167) | N13172);
assign N13170 = !N13167;
assign N13182 = !N11672;
assign N13174 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834;
assign N13166 = !(N13182 | N13174);
assign N13164 = !((N11667 | N13170) | N13166);
assign N13178 = !(N11500 & N11506);
assign x[22] = !(((N13181 | N13164) | N13151) & N13178);
assign N13152 = !N13151;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896 | a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834) ^ N11672;
assign x[21] = (N13154 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38]) | ((!N13154) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899) ^ N11677;
assign x[20] = (N13156 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37]) | ((!N13156) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608) ^ N11682;
assign x[19] = (N13155 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36]) | ((!N13155) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588) ^ N11687;
assign x[18] = (N13153 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35]) | ((!N13153) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831) ^ N11692;
assign x[17] = (N13154 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34]) | ((!N13154) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736) ^ N11697;
assign x[16] = (N13153 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33]) | ((!N13153) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911) ^ N11702;
assign x[15] = (N13155 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32]) | ((!N13155) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728) ^ N11707;
assign x[14] = (N13155 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31]) | ((!N13155) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820) ^ N11712;
assign x[13] = (N13154 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30]) | ((!N13154) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567) ^ N11717;
assign x[12] = (N13152 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29]) | ((!N13152) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579) ^ N11722;
assign x[11] = (N13152 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28]) | ((!N13152) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623;
assign x[10] = (N13152 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27]) | ((!N13152) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972;
assign x[9] = (N13154 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26]) | ((!N13154) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704;
assign x[8] = (N13156 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25]) | ((!N13156) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430;
assign x[7] = (N13155 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24]) | ((!N13155) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782;
assign x[6] = (N13153 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23]) | ((!N13153) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515;
assign x[5] = (N13153 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22]) | ((!N13153) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858;
assign x[4] = (N13153 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21]) | ((!N13153) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593;
assign x[3] = (N13155 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20]) | ((!N13155) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940;
assign x[2] = (N13156 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19]) | ((!N13156) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668;
assign x[1] = (N13154 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18]) | ((!N13154) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017;
assign x[0] = (N13152 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17]) | ((!N13152) & N13150);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | (!a_sign));
reg x_reg_23__I2278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__I2278_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23];
	end
assign x[23] = x_reg_23__I2278_QOUT;
reg x_reg_24__I2279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__I2279_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24];
	end
assign x[24] = x_reg_24__I2279_QOUT;
reg x_reg_25__I2280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_25__I2280_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25];
	end
assign x[25] = x_reg_25__I2280_QOUT;
reg x_reg_26__I2281_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__I2281_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26];
	end
assign x[26] = x_reg_26__I2281_QOUT;
reg x_reg_27__I2282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__I2282_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27];
	end
assign x[27] = x_reg_27__I2282_QOUT;
reg x_reg_28__I2283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__I2283_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28];
	end
assign x[28] = x_reg_28__I2283_QOUT;
reg x_reg_29__I2284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__I2284_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29];
	end
assign x[29] = x_reg_29__I2284_QOUT;
reg x_reg_30__I2285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I2285_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30];
	end
assign x[30] = x_reg_30__I2285_QOUT;
reg x_reg_31__I2286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I2286_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31];
	end
assign x[31] = x_reg_31__I2286_QOUT;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[0] = x[0];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[1] = x[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[2] = x[2];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[3] = x[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[4] = x[4];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[5] = x[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[6] = x[6];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[7] = x[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[8] = x[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[9] = x[9];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[10] = x[10];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[11] = x[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[12] = x[12];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[13] = x[13];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[14] = x[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[15] = x[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[19] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[20] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[24] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[39] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  vLTxTAvcrR8= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



