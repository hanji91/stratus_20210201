/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:10 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_4_0 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N446,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N448,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N455,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2353,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2384,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2393,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2402,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2404,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2516,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2518,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2576,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2578,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2581,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2584,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2585,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2586,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2587,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2588,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2590,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2591,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2593,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2595,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2597,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2599,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2600,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2602,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2604,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2608,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2609,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2611,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2614,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2615,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2616,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2617,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2619,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2620,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2621,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2623,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2624,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2626,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2628,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2629,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2630,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2632,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2633,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2635,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2636,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2638,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2641,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2642,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2643,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2644,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2647,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2649,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2650,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2655,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2656,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2659,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2661,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2665,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2666,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2670,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2671,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2673,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2674,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2675,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2677,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2678,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2679,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2680,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2681,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2682,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2683,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2684,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2685,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2686,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2688,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2689,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2691,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2694,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2695,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2696,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2699,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2701,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2702,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2704,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2706,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2708,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2709,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2711,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2712,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2713,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2714,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2715,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2717,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2719,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2720,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2721,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2724,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2726,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2727,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2731,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2732,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2735,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2744,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2745,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2747,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2749,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2752,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2754,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2759,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2761,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2771,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2774,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2778,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2781,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2782,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2784,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2786,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2788,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2793,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2797,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2801,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2802,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2803,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2805,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2807,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2815,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2817,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2818,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2820,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2821,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2824,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2826,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2829,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2830,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2832,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2833,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2837,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2838,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2842,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2843,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2844,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2845,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2855,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2858,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2860,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2862,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2864,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2867,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2869,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2874,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2877,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2879,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2880,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2883,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2885,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2891,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2894,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3203,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3204,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3205,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3206,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3208,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3211,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3212,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3213,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3214,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3216,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3217,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3218,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3219,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3222,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3224,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3226,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3229,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3230,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3231,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3232,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3234,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3235,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3236,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3238,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3239,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3242,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3243,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3245,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3251,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3252,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3253,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3255,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3257,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3259,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3260,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3262,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3263,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3264,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3265,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3266,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3268,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3269,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3270,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3271,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3272,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3273,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3274,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3275,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3276,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3278,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3279,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3280,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3281,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3282,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3283,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3285,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3286,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3287,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3288,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3290,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3291,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3293,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3294,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3298,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3301,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3302,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3303,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3304,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3305,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3306,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3309,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3310,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3311,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3312,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3314,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3316,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3318,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3321,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3322,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3323,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3325,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3327,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3329,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3331,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3332,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3334,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3336,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3339,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3340,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3341,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3343,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3346,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3347,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3348,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3352,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3353,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3354,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3356,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3357,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3358,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3359,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3360,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3361,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3362,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3363,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3364,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3365,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3368,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3369,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3370,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3371,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3372,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3374,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3375,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3377,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3379,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3380,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3383,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3385,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3386,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3390,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3391,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3396,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3398,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3401,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3405,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3406,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3407,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3415,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3420,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3423,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3431,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3435,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3436,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3443,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3447,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3465,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3469,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3470,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3472,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3476,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3490,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3497,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3505,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3509,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3513,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3516,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3519,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3522,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3527,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3531,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3539,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3543,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3544,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3551,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3554,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3557,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3561,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3566,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3567,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3572,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3575,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3576,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3585,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3586,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3587,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3591,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3595,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3604,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3607,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3610,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3614,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3615,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3630,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3635,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3644,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3645,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3650,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3651,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3652,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3654,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3655,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3659,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3660,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3667,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3677,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3678,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3688,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3689,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3693,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3697,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3698,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3701,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3707,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3711,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3727,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3732,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3736,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3738,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3740,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3746,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3747,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3748,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3755,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3764,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3774,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3780,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3781,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3782,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3784,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3786,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3788,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3794,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3797,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3799,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3801,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3802,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3803,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3804,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3805,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3807,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3810,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3813,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3816,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3817,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3818,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3820,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3821,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3822,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3824,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3826,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3830,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3832,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3833,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3834,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3835,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3837,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3840,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3842,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3843,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3844,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3845,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3847,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3856,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3859,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3860,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3862,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3866,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3869,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3873,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3876,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3877,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3879,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3880,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3882,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3883,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3884,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3885,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3890,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3892,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3894,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3896,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3899,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3900,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3901,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3902,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3903,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3904,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3905,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3906,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3907,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3909,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3912,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3913,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3915,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3916,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3917,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3918,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3919,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3920,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3922,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3923,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3924,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3925,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3928,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3929,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3930,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3933,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3934,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3935,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3936,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3937,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3939,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3940,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3941,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3942,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3943,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3944,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3945,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3946,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3949,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3950,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3951,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3953,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3954,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3957,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3959,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3962,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3963,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3964,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3965,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3966,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3968,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3969,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3970,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3971,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3972,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3973,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3975,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3976,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3977,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3979,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3980,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3981,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3982,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3984,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3985,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3986,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3988,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3989,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3992,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3994,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3995,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3996,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3997,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3998,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3999,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4000,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4002,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4004,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4005,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4006,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4007,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4008,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4009,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4010,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4011,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4012,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4015,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4016,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4017,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4018,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4019,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4020,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4021,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4022,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4025,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4027,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4028,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4029,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4030,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4031,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4032,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4033,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4035,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4036,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4037,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4038,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4039,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4041,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4043,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4046,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4047,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4048,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4049,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4050,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4051,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4053,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4055,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4057,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4059,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4060,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4061,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4062,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4066,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4067,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4068,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4070,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4073,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4074,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4075,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4076,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4079,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4080,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4082,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4083,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4084,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4085,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4086,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4087,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4088,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4090,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4091,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4092,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4093,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4094,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4095,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4096,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4098,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4101,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4102,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4103,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4104,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4107,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4108,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4109,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4110,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4111,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4113,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4114,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4116,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4117,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4120,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4121,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4122,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4123,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4124,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4125,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4126,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4127,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4128,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4130,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4131,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4133,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4134,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5062,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5067,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5070,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5076,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5084,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5092,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5095,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5098,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5102,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5105,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5111,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5114,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5119,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5126,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5130,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5135,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5138,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5144,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5151,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5154,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5155,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5161,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5162,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5165,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5166,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5167,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5169,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5171,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5172,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5173,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5175,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5176,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5177,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5178,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5179,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5182,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5183,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5184,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5185,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5187,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5189,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5190,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5192,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5193,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5194,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5195,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5196,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5197,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5198,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5199,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5201,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5203,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5204,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5206,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5207,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5208,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5209,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5211,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5212,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5214,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5215,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5216,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5217,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5218,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5220,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5221,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5223,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5224,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5226,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5228,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5229,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5231,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5232,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5233,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5235,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5236,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5237,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5238,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5240,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5241,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5242,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5244,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5245,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5247,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5248,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5249,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5250,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5252,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5254,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5255,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5256,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5257,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5258,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5260,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5261,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5263,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5264,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5265,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5266,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5267,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5268,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5269,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5270,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5272,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5273,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5274,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5276,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5277,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5279,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5280,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5281,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5283,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5284,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5286,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5287,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5289,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5290,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5291,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5293,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5295,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5296,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5297,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5299,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5300,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5301,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5302,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5303,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5304,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5305,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5307,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5308,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5309,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5310,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5311,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5312,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5313,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5315,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5316,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5318,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5319,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5320,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5321,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5323,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5324,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5325,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5326,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5327,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5328,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5330,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5332,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5333,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5335,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5337,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5338,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5339,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5340,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5341,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5342,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5343,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5344,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5345,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5346,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5347,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5349,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5352,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5353,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5354,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5356,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5357,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5358,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5361,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5362,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5363,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5364,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5366,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5367,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5368,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5370,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5371,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5372,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5374,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5377,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5379,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5382,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5384,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5385,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5386,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5388,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5390,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5391,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5393,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5396,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5398,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5399,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5400,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5401,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5721,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5724,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5726,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5728,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5729,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5731,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5732,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5735,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5736,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5738,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5739,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5740,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5743,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5744,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5745,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5747,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5748,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5749,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5751,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5752,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5754,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5756,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5758,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5760,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5764,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5766,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5771,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5772,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5774,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5777,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5778,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5780,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5782,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5784,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5785,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5788,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5792,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5793,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5795,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5797,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5799,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5801,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5802,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5804,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5805,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5807,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5810,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5813,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5816,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5818,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5820,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5821,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5822,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5824,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5825,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5829,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5832,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5833,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5834,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5836,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5837,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5838,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5840,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5841,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5842,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5844,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5845,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5847,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5849,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5855,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5856,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5858,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5859,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5862,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5863,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5864,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5867,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5870,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5872,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5873,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5874,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5875,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5877,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5879,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5880,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5882,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5883,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5884,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5885,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5888,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5889,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5890,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5892,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5894,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5896,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5897,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5898,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5899,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5901,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5902,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5903,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5904,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5905,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5906,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5909,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5910,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5912,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5913,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5914,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5915,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5916,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5917,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5918,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5919,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5920,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5921,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5922,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5925,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5926,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5927,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5928,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5929,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5930,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5931,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5932,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5933,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5935,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5936,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5937,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5938,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5939,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5941,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5942,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5944,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5946,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5947,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5948,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5949,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5950,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5952,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5953,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5954,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5955,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5956,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5958,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5959,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5960,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5961,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5962,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5963,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5964,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5965,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5966,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5967,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5968,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5969,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5970,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5971,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5974,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5975,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5976,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5977,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5978,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5979,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5980,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5981,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5982,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5983,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5984,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5985,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5986,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5987,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5988,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5991,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5992,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5993,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5994,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5995,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5996,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5997,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5998,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5999,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6000,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6001,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6002,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6003,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6005,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6007,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6008,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6009,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6010,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6011,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6012,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6014,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6015,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6016,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6017,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6019,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6020,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6021,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6022,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6024,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6025,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6026,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6027,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6028,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6029,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6030,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6031,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6032,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6034,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6035,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6036,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6037,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6038,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6039,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6040,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6041,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6044,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6045,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6046,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6047,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6049,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6050,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6051,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6053,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6054,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6055,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6056,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6058,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6059,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6060,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6061,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6062,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6063,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6064,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6065,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6067,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6068,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6069,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6070,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6071,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6072,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6073,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6074,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6076,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6077,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6078,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6079,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6080,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6082,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6083,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6084,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6085,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6086,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6087,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6089,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6090,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6091,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6093,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6094,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6095,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6096,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6098,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6099,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6100,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6101,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6102,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6103,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6104,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6105,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6107,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6109,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6110,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6113,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6114,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6115,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6116,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6117,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6118,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6119,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6121,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6122,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6124,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6125,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6126,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6128,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6129,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6130,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6131,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6132,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6134,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6135,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6136,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6137,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6138,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6139,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6140,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6141,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6143,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6144,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6145,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6146,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6147,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6148,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6149,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6150,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6151,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6152,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6153,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6154,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6155,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6156,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6158,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6159,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6160,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6161,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6162,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6163,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6165,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6167,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6168,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6169,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6170,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6171,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6172,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6175,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6177,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6178,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6180,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6186,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6187,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6193,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6194,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6202,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6207,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6210,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6212,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6221,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6231,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6237,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6238,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6240,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6241,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6248,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6250,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6254,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6261,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6263,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6271,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6274,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6279,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6280,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6282,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6288,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6292,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6293,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6294,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6300,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6313,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6314,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6319,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6322,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6323,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6325,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6330,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6335,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6336,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6338,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6340,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6343,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6346,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6351,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6352,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6356,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6364,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6368,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6375,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6377,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6384,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6385,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6388,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6398,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6399,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6402,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6406,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6410,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6411,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6418,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6423,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6426,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6431,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6439,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6440,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6443,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6448,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6460,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6461,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6462,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6463,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6466,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6470,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6471,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6472,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6485,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6499,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6506,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6507,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6510,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6515,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6516,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6517,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6519,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6520,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6521,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6522,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6524,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6525,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6527,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6528,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6529,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6530,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6532,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6533,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6534,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6535,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6536,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6537,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6538,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6540,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6541,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6543,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6544,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6545,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6546,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6547,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6549,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6550,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6551,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6552,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6553,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6555,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6556,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6557,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6558,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6559,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6560,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6561,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6562,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6563,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6564,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6565,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6566,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6569,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6570,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6572,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6573,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6574,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6575,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6577,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6578,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7414,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7416,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7423,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7427,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7436,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7445,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7461,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7505,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7512,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7525,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7528,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7548,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7549,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7552,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7556,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7561,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7566,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7602,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7607,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7609,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7624,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7625,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7631,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7636,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7637,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7642,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7647,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7656,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7662,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7663,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7665,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7673,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7676,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7688,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7692,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7694,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7696,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7698,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7709,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7711,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7713,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7716,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7720,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7739,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7758,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7778,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7785,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7786,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7795,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7804,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7825,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7843,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7859,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7860,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7873,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7876,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7889,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7902,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7903,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7909,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7921,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7922,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7924,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7925,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7926,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7927,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7929,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7940,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7943,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7946,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7949,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7959,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7961,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7962,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7963,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7967,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7969,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7970,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7972,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7979,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7980,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7984,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7987,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7988,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7990,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7993,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7996,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7997,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8001,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8004,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11575,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22792,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796;
wire N5603,N5608,N5613,N5618,N5623,N5628,N5633 
	,N5638,N5643,N11736,N11738,N11899,N11904,N11909,N11914 
	,N11919,N11924,N11929,N12012,N12014,N12065,N12067,N12072 
	,N12077,N12082,N12087,N12092,N12095,N12097,N12110,N12112 
	,N12118,N12120,N12136,N12138,N12144,N12146,N12154,N12156 
	,N12166,N12168,N12176,N12178,N12184,N12186,N12194,N12196 
	,N12206,N12268,N12270,N12272,N12294,N12298,N12320,N12354 
	,N12356,N12386,N12388,N12418,N12450,N12460,N12464,N12466 
	,N12538,N12586,N12599,N12605,N12607,N12609,N12647,N12669 
	,N12671,N12673,N12731,N12744,N12746,N12748,N12753,N12807 
	,N12823,N12825,N12827,N12885,N12893,N12895,N12897,N12963 
	,N13000,N13002,N13004,N13074,N13081,N13087,N13089,N13091 
	,N13094,N13104,N13189,N13197,N13199,N13201,N13205,N13207 
	,N13209,N13218,N13220,N13222,N13225,N13227,N13305,N13311 
	,N13319,N13335,N13337,N13424,N13430,N13432,N13436,N13448 
	,N13458,N13460,N13462,N13466,N13500,N13523,N13541,N13549 
	,N13551,N13555,N13557,N13583,N13585,N13587,N13591,N13593 
	,N13599,N13601,N13607,N13609,N13611,N13630,N13647,N13649 
	,N13659,N13673,N13675,N13681,N13685,N13689,N13693,N13697 
	,N13699,N13709,N13712,N13718,N13720,N13722,N13725,N13731 
	,N13733,N13735,N13761,N13763,N13769,N13771,N13773,N13777 
	,N13779,N13785,N13787,N13789,N13798,N13800,N13802,N13806 
	,N13808,N13810,N13822,N13824,N13835,N13837,N13842,N13852 
	,N13854,N13856,N13862,N13864,N13866,N13870,N13872,N13874 
	,N13878,N13880,N13882,N13888,N13890,N13892,N13896,N13898 
	,N13900,N14500,N14505,N14510,N14513,N14518,N14523,N14528 
	,N14533;
reg x_reg_L0_22__retimed_I7921_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7921_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355;
	end
assign N14533 = x_reg_L0_22__retimed_I7921_QOUT;
reg x_reg_L0_22__retimed_I7919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7919_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205;
	end
assign N14528 = x_reg_L0_22__retimed_I7919_QOUT;
reg x_reg_L0_22__retimed_I7917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7917_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132;
	end
assign N14523 = x_reg_L0_22__retimed_I7917_QOUT;
reg x_reg_L0_22__retimed_I7915_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7915_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397;
	end
assign N14518 = x_reg_L0_22__retimed_I7915_QOUT;
reg x_reg_L0_22__retimed_I7913_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7913_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164;
	end
assign N14513 = x_reg_L0_22__retimed_I7913_QOUT;
reg x_reg_L0_22__retimed_I7912_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7912_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219;
	end
assign N14510 = x_reg_L0_22__retimed_I7912_QOUT;
reg x_reg_L0_22__retimed_I7910_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7910_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365;
	end
assign N14505 = x_reg_L0_22__retimed_I7910_QOUT;
reg x_reg_L0_22__retimed_I7908_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7908_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292;
	end
assign N14500 = x_reg_L0_22__retimed_I7908_QOUT;
reg x_reg_L0_22__retimed_I7660_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7660_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[8];
	end
assign N13900 = x_reg_L0_22__retimed_I7660_QOUT;
reg x_reg_L0_22__retimed_I7659_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7659_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[8];
	end
assign N13898 = x_reg_L0_22__retimed_I7659_QOUT;
reg x_reg_L0_22__retimed_I7658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7658_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[8];
	end
assign N13896 = x_reg_L0_22__retimed_I7658_QOUT;
reg x_reg_L0_22__retimed_I7657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7657_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7949;
	end
assign N13892 = x_reg_L0_22__retimed_I7657_QOUT;
reg x_reg_L0_22__retimed_I7656_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7656_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[7];
	end
assign N13890 = x_reg_L0_22__retimed_I7656_QOUT;
reg x_reg_L0_22__retimed_I7655_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7655_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7445;
	end
assign N13888 = x_reg_L0_22__retimed_I7655_QOUT;
reg x_reg_L0_22__retimed_I7654_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7654_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5178;
	end
assign N13882 = x_reg_L0_22__retimed_I7654_QOUT;
reg x_reg_L0_22__retimed_I7653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7653_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5338;
	end
assign N13880 = x_reg_L0_22__retimed_I7653_QOUT;
reg x_reg_L0_22__retimed_I7652_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7652_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5371;
	end
assign N13878 = x_reg_L0_22__retimed_I7652_QOUT;
reg x_reg_L0_22__retimed_I7651_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7651_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5075;
	end
assign N13874 = x_reg_L0_22__retimed_I7651_QOUT;
reg x_reg_L0_22__retimed_I7650_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7650_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5264;
	end
assign N13872 = x_reg_L0_22__retimed_I7650_QOUT;
reg x_reg_L0_22__retimed_I7649_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7649_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5233;
	end
assign N13870 = x_reg_L0_22__retimed_I7649_QOUT;
reg x_reg_L0_22__retimed_I7648_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7648_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[9];
	end
assign N13866 = x_reg_L0_22__retimed_I7648_QOUT;
reg x_reg_L0_22__retimed_I7647_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7647_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[9];
	end
assign N13864 = x_reg_L0_22__retimed_I7647_QOUT;
reg x_reg_L0_22__retimed_I7646_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7646_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[9];
	end
assign N13862 = x_reg_L0_22__retimed_I7646_QOUT;
reg x_reg_L0_22__retimed_I7644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7644_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7789;
	end
assign N13856 = x_reg_L0_22__retimed_I7644_QOUT;
reg x_reg_L0_22__retimed_I7643_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7643_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7528;
	end
assign N13854 = x_reg_L0_22__retimed_I7643_QOUT;
reg x_reg_L0_22__retimed_I7642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7642_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7623;
	end
assign N13852 = x_reg_L0_22__retimed_I7642_QOUT;
reg x_reg_L0_22__retimed_I7638_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7638_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7925;
	end
assign N13842 = x_reg_L0_22__retimed_I7638_QOUT;
reg x_reg_L0_22__retimed_I7636_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7636_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7839;
	end
assign N13837 = x_reg_L0_22__retimed_I7636_QOUT;
reg x_reg_L0_22__retimed_I7635_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7635_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[8];
	end
assign N13835 = x_reg_L0_22__retimed_I7635_QOUT;
reg x_reg_L0_22__retimed_I7632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7632_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2588;
	end
assign N13824 = x_reg_L0_22__retimed_I7632_QOUT;
reg x_reg_L0_22__retimed_I7631_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7631_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2802;
	end
assign N13822 = x_reg_L0_22__retimed_I7631_QOUT;
reg x_reg_L0_22__retimed_I7630_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7630_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5236;
	end
assign N13810 = x_reg_L0_22__retimed_I7630_QOUT;
reg x_reg_L0_22__retimed_I7629_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7629_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5372;
	end
assign N13808 = x_reg_L0_22__retimed_I7629_QOUT;
reg x_reg_L0_22__retimed_I7628_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7628_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5166;
	end
assign N13806 = x_reg_L0_22__retimed_I7628_QOUT;
reg x_reg_L0_22__retimed_I7627_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7627_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5363;
	end
assign N13802 = x_reg_L0_22__retimed_I7627_QOUT;
reg x_reg_L0_22__retimed_I7626_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7626_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5158;
	end
assign N13800 = x_reg_L0_22__retimed_I7626_QOUT;
reg x_reg_L0_22__retimed_I7625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7625_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5291;
	end
assign N13798 = x_reg_L0_22__retimed_I7625_QOUT;
reg x_reg_L0_22__retimed_I7622_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7622_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5378;
	end
assign N13789 = x_reg_L0_22__retimed_I7622_QOUT;
reg x_reg_L0_22__retimed_I7621_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7621_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5304;
	end
assign N13787 = x_reg_L0_22__retimed_I7621_QOUT;
reg x_reg_L0_22__retimed_I7620_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7620_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5172;
	end
assign N13785 = x_reg_L0_22__retimed_I7620_QOUT;
reg x_reg_L0_22__retimed_I7618_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7618_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[10];
	end
assign N13779 = x_reg_L0_22__retimed_I7618_QOUT;
reg x_reg_L0_22__retimed_I7617_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7617_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[10];
	end
assign N13777 = x_reg_L0_22__retimed_I7617_QOUT;
reg x_reg_L0_22__retimed_I7616_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7616_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5388;
	end
assign N13773 = x_reg_L0_22__retimed_I7616_QOUT;
reg x_reg_L0_22__retimed_I7615_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7615_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5238;
	end
assign N13771 = x_reg_L0_22__retimed_I7615_QOUT;
reg x_reg_L0_22__retimed_I7614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7614_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5062;
	end
assign N13769 = x_reg_L0_22__retimed_I7614_QOUT;
reg x_reg_L0_22__retimed_I7612_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7612_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5327;
	end
assign N13763 = x_reg_L0_22__retimed_I7612_QOUT;
reg x_reg_L0_22__retimed_I7611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7611_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5151;
	end
assign N13761 = x_reg_L0_22__retimed_I7611_QOUT;
reg x_reg_L0_22__retimed_I7602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7602_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5844;
	end
assign N13735 = x_reg_L0_22__retimed_I7602_QOUT;
reg x_reg_L0_22__retimed_I7601_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7601_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6330;
	end
assign N13733 = x_reg_L0_22__retimed_I7601_QOUT;
reg x_reg_L0_22__retimed_I7600_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7600_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6206;
	end
assign N13731 = x_reg_L0_22__retimed_I7600_QOUT;
reg x_reg_L0_22__retimed_I7598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7598_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322;
	end
assign N13725 = x_reg_L0_22__retimed_I7598_QOUT;
reg x_reg_L0_22__retimed_I7597_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7597_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5112;
	end
assign N13722 = x_reg_L0_22__retimed_I7597_QOUT;
reg x_reg_L0_22__retimed_I7596_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7596_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5123;
	end
assign N13720 = x_reg_L0_22__retimed_I7596_QOUT;
reg x_reg_L0_22__retimed_I7595_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7595_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5313;
	end
assign N13718 = x_reg_L0_22__retimed_I7595_QOUT;
reg x_reg_L0_22__retimed_I7593_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7593_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246;
	end
assign N13712 = x_reg_L0_22__retimed_I7593_QOUT;
reg x_reg_L0_22__retimed_I7592_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7592_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5179;
	end
assign N13709 = x_reg_L0_22__retimed_I7592_QOUT;
reg x_reg_L0_22__retimed_I7588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7588_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5184;
	end
assign N13699 = x_reg_L0_22__retimed_I7588_QOUT;
reg x_reg_L0_22__retimed_I7587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7587_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5320;
	end
assign N13697 = x_reg_L0_22__retimed_I7587_QOUT;
reg x_reg_L0_22__retimed_I7586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7586_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5203;
	end
assign N13693 = x_reg_L0_22__retimed_I7586_QOUT;
reg x_reg_L0_22__retimed_I7584_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7584_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5395;
	end
assign N13689 = x_reg_L0_22__retimed_I7584_QOUT;
reg x_reg_L0_22__retimed_I7583_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7583_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5069;
	end
assign N13685 = x_reg_L0_22__retimed_I7583_QOUT;
reg x_reg_L0_22__retimed_I7581_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7581_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5269;
	end
assign N13681 = x_reg_L0_22__retimed_I7581_QOUT;
reg x_reg_L0_22__retimed_I7579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7579_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5144;
	end
assign N13675 = x_reg_L0_22__retimed_I7579_QOUT;
reg x_reg_L0_22__retimed_I7578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7578_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5130;
	end
assign N13673 = x_reg_L0_22__retimed_I7578_QOUT;
reg x_reg_L0_22__retimed_I7573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7573_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5150;
	end
assign N13659 = x_reg_L0_22__retimed_I7573_QOUT;
reg x_reg_L0_22__retimed_I7569_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7569_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[11];
	end
assign N13649 = x_reg_L0_22__retimed_I7569_QOUT;
reg x_reg_L0_22__retimed_I7568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7568_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[11];
	end
assign N13647 = x_reg_L0_22__retimed_I7568_QOUT;
reg x_reg_L0_22__retimed_I7561_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7561_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5197;
	end
assign N13630 = x_reg_L0_22__retimed_I7561_QOUT;
reg x_reg_L0_22__retimed_I7555_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7555_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6044;
	end
assign N13611 = x_reg_L0_22__retimed_I7555_QOUT;
reg x_reg_L0_22__retimed_I7554_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7554_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6030;
	end
assign N13609 = x_reg_L0_22__retimed_I7554_QOUT;
reg x_reg_L0_22__retimed_I7553_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7553_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6535;
	end
assign N13607 = x_reg_L0_22__retimed_I7553_QOUT;
reg x_reg_L0_22__retimed_I7551_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7551_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5198;
	end
assign N13601 = x_reg_L0_22__retimed_I7551_QOUT;
reg x_reg_L0_22__retimed_I7550_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7550_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5133;
	end
assign N13599 = x_reg_L0_22__retimed_I7550_QOUT;
reg x_reg_L0_22__retimed_I7548_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7548_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5122;
	end
assign N13593 = x_reg_L0_22__retimed_I7548_QOUT;
reg x_reg_L0_22__retimed_I7547_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7547_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5389;
	end
assign N13591 = x_reg_L0_22__retimed_I7547_QOUT;
reg x_reg_L0_22__retimed_I7546_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7546_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5762;
	end
assign N13587 = x_reg_L0_22__retimed_I7546_QOUT;
reg x_reg_L0_22__retimed_I7545_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7545_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6246;
	end
assign N13585 = x_reg_L0_22__retimed_I7545_QOUT;
reg x_reg_L0_22__retimed_I7544_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7544_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6231;
	end
assign N13583 = x_reg_L0_22__retimed_I7544_QOUT;
reg x_reg_L0_22__retimed_I7534_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7534_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5396;
	end
assign N13557 = x_reg_L0_22__retimed_I7534_QOUT;
reg x_reg_L0_22__retimed_I7533_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7533_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5260;
	end
assign N13555 = x_reg_L0_22__retimed_I7533_QOUT;
reg x_reg_L0_22__retimed_I7532_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7532_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5370;
	end
assign N13551 = x_reg_L0_22__retimed_I7532_QOUT;
reg x_reg_L0_22__retimed_I7531_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7531_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5223;
	end
assign N13549 = x_reg_L0_22__retimed_I7531_QOUT;
reg x_reg_L0_22__retimed_I7528_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7528_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5311;
	end
assign N13541 = x_reg_L0_22__retimed_I7528_QOUT;
reg x_reg_L0_22__retimed_I7521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7521_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5296;
	end
assign N13523 = x_reg_L0_22__retimed_I7521_QOUT;
reg x_reg_L0_22__retimed_I7512_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7512_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[12];
	end
assign N13500 = x_reg_L0_22__retimed_I7512_QOUT;
reg x_reg_L0_22__retimed_I7500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7500_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N477;
	end
assign N13466 = x_reg_L0_22__retimed_I7500_QOUT;
reg x_reg_L0_22__retimed_I7499_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7499_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6228;
	end
assign N13462 = x_reg_L0_22__retimed_I7499_QOUT;
reg x_reg_L0_22__retimed_I7498_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7498_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5950;
	end
assign N13460 = x_reg_L0_22__retimed_I7498_QOUT;
reg x_reg_L0_22__retimed_I7497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7497_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5853;
	end
assign N13458 = x_reg_L0_22__retimed_I7497_QOUT;
reg x_reg_L0_22__retimed_I7494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7494_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5148;
	end
assign N13448 = x_reg_L0_22__retimed_I7494_QOUT;
reg x_reg_L0_22__retimed_I7489_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7489_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5139;
	end
assign N13436 = x_reg_L0_22__retimed_I7489_QOUT;
reg x_reg_L0_22__retimed_I7488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7488_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5387;
	end
assign N13432 = x_reg_L0_22__retimed_I7488_QOUT;
reg x_reg_L0_22__retimed_I7487_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7487_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5143;
	end
assign N13430 = x_reg_L0_22__retimed_I7487_QOUT;
reg x_reg_L0_22__retimed_I7485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7485_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5215;
	end
assign N13424 = x_reg_L0_22__retimed_I7485_QOUT;
reg x_reg_L0_22__retimed_I7452_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7452_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5087;
	end
assign N13337 = x_reg_L0_22__retimed_I7452_QOUT;
reg x_reg_L0_22__retimed_I7451_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7451_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5157;
	end
assign N13335 = x_reg_L0_22__retimed_I7451_QOUT;
reg x_reg_L0_22__retimed_I7445_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7445_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5361;
	end
assign N13319 = x_reg_L0_22__retimed_I7445_QOUT;
reg x_reg_L0_22__retimed_I7442_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7442_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5381;
	end
assign N13311 = x_reg_L0_22__retimed_I7442_QOUT;
reg x_reg_L0_22__retimed_I7440_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7440_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5305;
	end
assign N13305 = x_reg_L0_22__retimed_I7440_QOUT;
reg x_reg_L1_16__retimed_I7411_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I7411_QOUT <= N11929;
	end
assign N13227 = x_reg_L1_16__retimed_I7411_QOUT;
reg x_reg_L1_16__retimed_I7410_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I7410_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854;
	end
assign N13225 = x_reg_L1_16__retimed_I7410_QOUT;
reg x_reg_L0_22__retimed_I7409_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7409_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5235;
	end
assign N13222 = x_reg_L0_22__retimed_I7409_QOUT;
reg x_reg_L0_22__retimed_I7408_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7408_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5171;
	end
assign N13220 = x_reg_L0_22__retimed_I7408_QOUT;
reg x_reg_L0_22__retimed_I7407_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7407_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5303;
	end
assign N13218 = x_reg_L0_22__retimed_I7407_QOUT;
reg x_reg_L0_22__retimed_I7404_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7404_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6325;
	end
assign N13209 = x_reg_L0_22__retimed_I7404_QOUT;
reg x_reg_L0_22__retimed_I7403_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7403_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6418;
	end
assign N13207 = x_reg_L0_22__retimed_I7403_QOUT;
reg x_reg_L0_22__retimed_I7402_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7402_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5948;
	end
assign N13205 = x_reg_L0_22__retimed_I7402_QOUT;
reg x_reg_L0_22__retimed_I7401_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7401_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6413;
	end
assign N13201 = x_reg_L0_22__retimed_I7401_QOUT;
reg x_reg_L0_22__retimed_I7400_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7400_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6514;
	end
assign N13199 = x_reg_L0_22__retimed_I7400_QOUT;
reg x_reg_L0_22__retimed_I7399_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7399_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6035;
	end
assign N13197 = x_reg_L0_22__retimed_I7399_QOUT;
reg x_reg_L0_22__retimed_I7396_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7396_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5104;
	end
assign N13189 = x_reg_L0_22__retimed_I7396_QOUT;
reg x_reg_L0_22__retimed_I7364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7364_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086;
	end
assign N13104 = x_reg_L0_22__retimed_I7364_QOUT;
reg x_reg_L0_22__retimed_I7360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7360_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N478;
	end
assign N13094 = x_reg_L0_22__retimed_I7360_QOUT;
reg x_reg_L0_22__retimed_I7359_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7359_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6021;
	end
assign N13091 = x_reg_L0_22__retimed_I7359_QOUT;
reg x_reg_L0_22__retimed_I7358_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7358_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5739;
	end
assign N13089 = x_reg_L0_22__retimed_I7358_QOUT;
reg x_reg_L0_22__retimed_I7357_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7357_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6509;
	end
assign N13087 = x_reg_L0_22__retimed_I7357_QOUT;
reg x_reg_L0_22__retimed_I7355_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7355_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278;
	end
assign N13081 = x_reg_L0_22__retimed_I7355_QOUT;
reg x_reg_L0_22__retimed_I7352_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7352_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N479;
	end
assign N13074 = x_reg_L0_22__retimed_I7352_QOUT;
reg x_reg_L0_22__retimed_I7327_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7327_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6110;
	end
assign N13004 = x_reg_L0_22__retimed_I7327_QOUT;
reg x_reg_L0_22__retimed_I7326_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7326_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6209;
	end
assign N13002 = x_reg_L0_22__retimed_I7326_QOUT;
reg x_reg_L0_22__retimed_I7325_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7325_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5736;
	end
assign N13000 = x_reg_L0_22__retimed_I7325_QOUT;
reg x_reg_L0_22__retimed_I7311_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7311_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N480;
	end
assign N12963 = x_reg_L0_22__retimed_I7311_QOUT;
reg x_reg_L0_22__retimed_I7287_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7287_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5831;
	end
assign N12897 = x_reg_L0_22__retimed_I7287_QOUT;
reg x_reg_L0_22__retimed_I7286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7286_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6297;
	end
assign N12895 = x_reg_L0_22__retimed_I7286_QOUT;
reg x_reg_L0_22__retimed_I7285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7285_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6315;
	end
assign N12893 = x_reg_L0_22__retimed_I7285_QOUT;
reg x_reg_L0_22__retimed_I7282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7282_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N481;
	end
assign N12885 = x_reg_L0_22__retimed_I7282_QOUT;
reg x_reg_L0_22__retimed_I7261_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7261_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6029;
	end
assign N12827 = x_reg_L0_22__retimed_I7261_QOUT;
reg x_reg_L0_22__retimed_I7260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7260_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6017;
	end
assign N12825 = x_reg_L0_22__retimed_I7260_QOUT;
reg x_reg_L0_22__retimed_I7259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7259_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6517;
	end
assign N12823 = x_reg_L0_22__retimed_I7259_QOUT;
reg x_reg_L0_22__retimed_I7253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7253_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N482;
	end
assign N12807 = x_reg_L0_22__retimed_I7253_QOUT;
reg x_reg_L0_22__retimed_I7234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7234_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5101;
	end
assign N12753 = x_reg_L0_22__retimed_I7234_QOUT;
reg x_reg_L0_22__retimed_I7232_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7232_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5855;
	end
assign N12748 = x_reg_L0_22__retimed_I7232_QOUT;
reg x_reg_L0_22__retimed_I7231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7231_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6218;
	end
assign N12746 = x_reg_L0_22__retimed_I7231_QOUT;
reg x_reg_L0_22__retimed_I7230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7230_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6343;
	end
assign N12744 = x_reg_L0_22__retimed_I7230_QOUT;
reg x_reg_L0_22__retimed_I7225_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7225_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N483;
	end
assign N12731 = x_reg_L0_22__retimed_I7225_QOUT;
reg x_reg_L0_22__retimed_I7205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7205_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6167;
	end
assign N12673 = x_reg_L0_22__retimed_I7205_QOUT;
reg x_reg_L0_22__retimed_I7204_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7204_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6041;
	end
assign N12671 = x_reg_L0_22__retimed_I7204_QOUT;
reg x_reg_L0_22__retimed_I7203_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7203_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5792;
	end
assign N12669 = x_reg_L0_22__retimed_I7203_QOUT;
reg x_reg_L0_22__retimed_I7195_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7195_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N484;
	end
assign N12647 = x_reg_L0_22__retimed_I7195_QOUT;
reg x_reg_L0_22__retimed_I7182_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7182_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6103;
	end
assign N12609 = x_reg_L0_22__retimed_I7182_QOUT;
reg x_reg_L0_22__retimed_I7181_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7181_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6358;
	end
assign N12607 = x_reg_L0_22__retimed_I7181_QOUT;
reg x_reg_L0_22__retimed_I7180_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7180_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5732;
	end
assign N12605 = x_reg_L0_22__retimed_I7180_QOUT;
reg x_reg_L0_22__retimed_I7178_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7178_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234;
	end
assign N12599 = x_reg_L0_22__retimed_I7178_QOUT;
reg x_reg_L0_22__retimed_I7173_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7173_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N485;
	end
assign N12586 = x_reg_L0_22__retimed_I7173_QOUT;
reg x_reg_L0_22__retimed_I7156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7156_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N486;
	end
assign N12538 = x_reg_L0_22__retimed_I7156_QOUT;
reg x_reg_L0_22__retimed_I7131_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7131_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[26];
	end
assign N12466 = x_reg_L0_22__retimed_I7131_QOUT;
reg x_reg_L0_22__retimed_I7130_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7130_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[26];
	end
assign N12464 = x_reg_L0_22__retimed_I7130_QOUT;
reg x_reg_L0_22__retimed_I7129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7129_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[25];
	end
assign N12460 = x_reg_L0_22__retimed_I7129_QOUT;
reg x_reg_L0_22__retimed_I7125_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7125_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N487;
	end
assign N12450 = x_reg_L0_22__retimed_I7125_QOUT;
reg x_reg_L0_22__retimed_I7114_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7114_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N488;
	end
assign N12418 = x_reg_L0_22__retimed_I7114_QOUT;
reg x_reg_L0_22__retimed_I7104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7104_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7416;
	end
assign N12388 = x_reg_L0_22__retimed_I7104_QOUT;
reg x_reg_L0_22__retimed_I7103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7103_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N489;
	end
assign N12386 = x_reg_L0_22__retimed_I7103_QOUT;
reg x_reg_L0_22__retimed_I7093_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7093_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7946;
	end
assign N12356 = x_reg_L0_22__retimed_I7093_QOUT;
reg x_reg_L0_22__retimed_I7092_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7092_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N490;
	end
assign N12354 = x_reg_L0_22__retimed_I7092_QOUT;
reg x_reg_L0_22__retimed_I7080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7080_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7548;
	end
assign N12320 = x_reg_L0_22__retimed_I7080_QOUT;
reg x_reg_L0_22__retimed_I7073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7073_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7570;
	end
assign N12298 = x_reg_L0_22__retimed_I7073_QOUT;
reg x_reg_L0_22__retimed_I7071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7071_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7474;
	end
assign N12294 = x_reg_L0_22__retimed_I7071_QOUT;
reg x_reg_L0_22__retimed_I7064_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7064_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7478;
	end
assign N12272 = x_reg_L0_22__retimed_I7064_QOUT;
reg x_reg_L0_22__retimed_I7063_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7063_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7479;
	end
assign N12270 = x_reg_L0_22__retimed_I7063_QOUT;
reg x_reg_L0_22__retimed_I7062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7062_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7996;
	end
assign N12268 = x_reg_L0_22__retimed_I7062_QOUT;
reg x_reg_L0_22__retimed_I7040_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7040_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8001;
	end
assign N12206 = x_reg_L0_22__retimed_I7040_QOUT;
reg x_reg_L0_22__retimed_I7036_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7036_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7532;
	end
assign N12196 = x_reg_L0_22__retimed_I7036_QOUT;
reg x_reg_L0_22__retimed_I7035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7035_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7798;
	end
assign N12194 = x_reg_L0_22__retimed_I7035_QOUT;
reg x_reg_L1_22__retimed_I7032_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7032_QOUT <= N12156;
	end
assign N12186 = x_reg_L1_22__retimed_I7032_QOUT;
reg x_reg_L1_22__retimed_I7031_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7031_QOUT <= N12154;
	end
assign N12184 = x_reg_L1_22__retimed_I7031_QOUT;
reg x_reg_L0_22__retimed_I7029_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7029_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931;
	end
assign N12178 = x_reg_L0_22__retimed_I7029_QOUT;
reg x_reg_L0_22__retimed_I7028_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7028_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581;
	end
assign N12176 = x_reg_L0_22__retimed_I7028_QOUT;
reg x_reg_L1_22__retimed_I7025_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7025_QOUT <= N12138;
	end
assign N12168 = x_reg_L1_22__retimed_I7025_QOUT;
reg x_reg_L1_22__retimed_I7024_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7024_QOUT <= N12136;
	end
assign N12166 = x_reg_L1_22__retimed_I7024_QOUT;
reg x_reg_L0_22__retimed_I7020_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7020_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722;
	end
assign N12156 = x_reg_L0_22__retimed_I7020_QOUT;
reg x_reg_L0_22__retimed_I7019_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7019_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982;
	end
assign N12154 = x_reg_L0_22__retimed_I7019_QOUT;
reg x_reg_L1_22__retimed_I7016_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7016_QOUT <= N12120;
	end
assign N12146 = x_reg_L1_22__retimed_I7016_QOUT;
reg x_reg_L1_22__retimed_I7015_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7015_QOUT <= N12118;
	end
assign N12144 = x_reg_L1_22__retimed_I7015_QOUT;
reg x_reg_L0_22__retimed_I7013_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7013_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514;
	end
assign N12138 = x_reg_L0_22__retimed_I7013_QOUT;
reg x_reg_L0_22__retimed_I7012_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7012_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775;
	end
assign N12136 = x_reg_L0_22__retimed_I7012_QOUT;
reg x_reg_L0_22__retimed_I7006_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7006_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484;
	end
assign N12120 = x_reg_L0_22__retimed_I7006_QOUT;
reg x_reg_L0_22__retimed_I7005_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7005_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911;
	end
assign N12118 = x_reg_L0_22__retimed_I7005_QOUT;
reg x_reg_L1_22__retimed_I7003_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7003_QOUT <= N12067;
	end
assign N12112 = x_reg_L1_22__retimed_I7003_QOUT;
reg x_reg_L1_22__retimed_I7002_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7002_QOUT <= N12065;
	end
assign N12110 = x_reg_L1_22__retimed_I7002_QOUT;
reg x_reg_L1_17__retimed_I6997_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I6997_QOUT <= N11924;
	end
assign N12097 = x_reg_L1_17__retimed_I6997_QOUT;
reg x_reg_L1_17__retimed_I6996_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I6996_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7692;
	end
assign N12095 = x_reg_L1_17__retimed_I6996_QOUT;
reg x_reg_L1_18__retimed_I6995_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I6995_QOUT <= N11919;
	end
assign N12092 = x_reg_L1_18__retimed_I6995_QOUT;
reg x_reg_L1_19__retimed_I6993_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I6993_QOUT <= N11914;
	end
assign N12087 = x_reg_L1_19__retimed_I6993_QOUT;
reg x_reg_L1_20__retimed_I6991_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I6991_QOUT <= N11909;
	end
assign N12082 = x_reg_L1_20__retimed_I6991_QOUT;
reg x_reg_L1_21__retimed_I6989_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I6989_QOUT <= N11904;
	end
assign N12077 = x_reg_L1_21__retimed_I6989_QOUT;
reg x_reg_L1_22__retimed_I6987_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I6987_QOUT <= N11899;
	end
assign N12072 = x_reg_L1_22__retimed_I6987_QOUT;
reg x_reg_L0_22__retimed_I6985_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6985_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755;
	end
assign N12067 = x_reg_L0_22__retimed_I6985_QOUT;
reg x_reg_L0_22__retimed_I6984_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6984_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491;
	end
assign N12065 = x_reg_L0_22__retimed_I6984_QOUT;
reg x_reg_L1_22__retimed_I6962_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I6962_QOUT <= N11738;
	end
assign N12014 = x_reg_L1_22__retimed_I6962_QOUT;
reg x_reg_L1_22__retimed_I6961_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I6961_QOUT <= N11736;
	end
assign N12012 = x_reg_L1_22__retimed_I6961_QOUT;
reg x_reg_L0_16__retimed_I6928_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I6928_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7993;
	end
assign N11929 = x_reg_L0_16__retimed_I6928_QOUT;
reg x_reg_L0_17__retimed_I6926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I6926_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7654;
	end
assign N11924 = x_reg_L0_17__retimed_I6926_QOUT;
reg x_reg_L0_18__retimed_I6924_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I6924_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7924;
	end
assign N11919 = x_reg_L0_18__retimed_I6924_QOUT;
reg x_reg_L0_19__retimed_I6922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I6922_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7572;
	end
assign N11914 = x_reg_L0_19__retimed_I6922_QOUT;
reg x_reg_L0_20__retimed_I6920_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I6920_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7962;
	end
assign N11909 = x_reg_L0_20__retimed_I6920_QOUT;
reg x_reg_L0_21__retimed_I6918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6918_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7505;
	end
assign N11904 = x_reg_L0_21__retimed_I6918_QOUT;
reg x_reg_L0_22__retimed_I6916_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6916_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7765;
	end
assign N11899 = x_reg_L0_22__retimed_I6916_QOUT;
reg x_reg_L0_22__retimed_I6847_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6847_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29;
	end
assign N11738 = x_reg_L0_22__retimed_I6847_QOUT;
reg x_reg_L0_22__retimed_I6846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6846_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__67;
	end
assign N11736 = x_reg_L0_22__retimed_I6846_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2353 = !(a_exp[7] & a_exp[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2355 = ((a_exp[4] & a_exp[3]) & a_exp[2]) & a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11575 = !((a_exp[6] & a_exp[5]) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2355);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2353 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11575);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2376 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2395 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2384 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2404 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2387 = !(((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2376 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2395) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2384) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2404);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2389 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2393 = !(((a_man[0] | a_man[1]) | a_man[2]) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2389);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 = !(a_man[18] | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2408 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2402 = !((((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381) | a_man[16]) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2408) | a_man[15]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2378 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2393 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2402);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0] = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2387 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2378);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0] | (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425 = !a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112 = !a_man[21];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409 = !a_man[20];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 = !a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 = !a_man[18];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 = !(a_man[17] | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 = !a_man[17];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 = !a_man[16];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3456 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4009 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3212 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3456 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4009 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 = !(a_man[16] & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3847 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3627 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3807 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3847 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3627 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3821 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3212 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3807 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4020 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3250 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4020 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (a_man[19] & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052 = !(a_man[19] | a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4010 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3413 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3250 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4010 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3821 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3413 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7825 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3666 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013 = !(a_man[17] & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3280 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3414 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3666 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3280 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3827 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4005 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3827 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4021 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3414 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4005 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3455 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3281 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3624 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3455 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3281 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4021 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3624 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7987 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7962} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7825} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7987};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3625 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3294 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3625 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3356 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3356 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3824 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3294 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3824 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7505 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[16]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3251 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3944 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3251 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3273 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3647 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3273 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3416 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3605 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3647 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3416 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3620 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3944 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3605 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3820 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3361 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3979 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3820 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3361 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3848 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3812 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3848 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3211 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3979 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3812 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3620 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3211 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3980 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 = !(a_man[17] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 = !((a_man[17] & a_man[16]) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3609 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3743 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3980 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3609 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3438 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3214 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3396 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3438 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3214 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3408 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3743 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3396 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3618 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4092 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3779 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3618 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4092 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3651 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3648 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3610 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3651 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3648 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3943 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3779 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3610 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N496 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3408 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3943 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7686} = {1'B0, 1'B1} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N496};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7572 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] = !a_man[15];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3375 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3398 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3539 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3375 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3398 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3233 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3946 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4131 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3233 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3946 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3208 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3539 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4131 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3406 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3885 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3574 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3406 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3885 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3443 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3439 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3399 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3443 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3439 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3742 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3574 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3399 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N495 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3208 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3742 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3587 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[17] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3587 & a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6466 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 = !a_man[14];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[17];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6059 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 = !a_man[13];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3527 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4117 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3604 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3527 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4117 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[16] = !(a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3604);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6085 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[16]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6524, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6335} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6059} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6085};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[33], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[32]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6466} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6524};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7696, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7556} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N495} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[33]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7848, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7785} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7556};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7696} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7848} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7686};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4108 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4133 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3335 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4108 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4133 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3966 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[18] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3930 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3966 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3942 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3335 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3930 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3205 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3686 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3374 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3205 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3686 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3236 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3234 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4134 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3236 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3234 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3538 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3374 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4134 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N494 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3942 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3538 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6520 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 = !a_man[12];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3561 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3321 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3561 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3913 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3394 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3321 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3913 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3846 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3526 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3846 | a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[15] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3394 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3526 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6577 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[15]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6255, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6068} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6520} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6577};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6114 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 = !a_man[11];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3359 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3917 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4047 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3359 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3917 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3748 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3708 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3748 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4130 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4047 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3708 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4090 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4120 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3320 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4090 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4120 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[14] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4130 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3320 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6198 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[14]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6480, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6289} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6114} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6198};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[16];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6547 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5771, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6446} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6547} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6480} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6068};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[32], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[31]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6255} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6335} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5771};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7770, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7634} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[32]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[32]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7453, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7887} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7634};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7770} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7453} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7785};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7654 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4123 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3900 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4123 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3933 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4061 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3900 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3933 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3765 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3862 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3727 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3765 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3862 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3740 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4061 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3727 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3937 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3478 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4107 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3937 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3478 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3968 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3934 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3968 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3334 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4107 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3934 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N493 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3740 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3334 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[15];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6171 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6141 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6574 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 = !a_man[10];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4091 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3713 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3843 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4091 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3713 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3506 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3928 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3843 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3506 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3723 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3985 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3883 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3985 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3918 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4046 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3883 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3918 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[13] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3928 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4046 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5823 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[13]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6324, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6135} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6574} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5823};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5993, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5805} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6141} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6171} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6324};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5766 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5738 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[14];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5796 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5838, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6512} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5738} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5766} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5796};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6369, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6180} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6289} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5838} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5805};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[31], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[30]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5993} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6446} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6369};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7843, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7716} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[31]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[31]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7665, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7980} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7716};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7798} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7843} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7665} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7887};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3329 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3698 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3329 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3729 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3860 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3698 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3729 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3557 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3663 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3523 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3557 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3663 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3537 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3860 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3523 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3293 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3738 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3293 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3271 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3899 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3738 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3271 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3767 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4087 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3730 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3767 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4087 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4060 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3899 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3730 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N492 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3537 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4060 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6168 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 = !a_man[9];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3884 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3510 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3644 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3884 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3510 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3340 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3298 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3340 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3725 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3644 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3298 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3521 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3786 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3684 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3521 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3786 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3982 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3714 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3982 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3842 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3684 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3714 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[12] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3725 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3842 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6308 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[12]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5790, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6463} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6168} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6308};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6223 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6196 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6250 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6163, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5978} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6196} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6223} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6250};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6212, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6026} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5790} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6135} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6163};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5763 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 = !a_man[8];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5793 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5742, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6416} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5763} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5793};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[13];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6279 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6544, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6356} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6279} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5742} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6463};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5729, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6403} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6512} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6544} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6026};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[30], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[29]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6212} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6180} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5729};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7927, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7791} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[30]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[30]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7878, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7478} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N492} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7791};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7532, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8001} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7927} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7878} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7980};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736 = (!N12194) ^ N12196;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3514 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3495 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3514 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3529 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3661 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3495 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3529 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3357 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3453 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3318 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3357 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3453 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3332 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3661 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3318 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3535 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4000 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3697 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3535 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4000 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3564 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3881 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3530 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3564 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3881 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3859 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3697 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3530 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N491 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3332 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3859 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5875 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6221 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 = !a_man[7];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3477 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4029 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3230 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3477 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4029 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3866 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3559 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3826 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3866 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3559 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3316 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3230 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3826 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4038 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3379 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3268 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4038 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3379 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3460 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3577 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3304 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3460 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3577 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3434 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3268 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3304 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[10] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3316 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3434 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6419 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[10]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6185, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5997} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6221} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6419};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[12];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5905 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6494, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6305} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5875} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5905};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5821 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3685 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3303 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3435 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3685 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3303 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4068 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3766 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4025 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4068 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3766 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3522 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3435 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4025 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3314 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3580 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3476 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3314 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3580 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3781 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[18] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3511 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3781 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3643 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3476 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3511 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[11] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3522 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3643 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5932 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[11]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5848 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6117, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5930} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5932} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5821} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5848};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6054, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5867} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6117} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5978};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6276 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6248 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6306 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6559, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6373} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6248} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6276} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6306};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6336 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5818 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 = !a_man[6];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3269 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3832 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3963 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3269 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3832 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3667 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3358 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3626 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3667 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3358 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4041 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3963 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3626 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3428 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4113 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3998 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3428 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4113 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3256 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3378 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4031 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3256 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3378 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3229 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3998 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4031 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[9] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4041 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3229 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6039 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[9]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6245, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6056} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5818} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6039};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6364 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6072, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5883} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6245} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6336} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6364};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6008, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5820} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6416} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6559} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6072};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6432, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6243} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6356} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6008} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5867};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[29], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[28]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6054} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6403} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6432};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7996, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7873} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[29]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[29]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7479, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7570} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N491} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7873};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605} = {1'B0, N12268} + {1'B0, N12270} + {1'B0, N12272};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3286 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3322 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3452 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3286 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3322 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3235 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4086 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3235 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3247 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4043 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4086 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3247 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4059 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3452 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4043 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3328 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3253 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3803 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3253 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3494 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3328 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3803 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3703 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3363 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3703 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3682 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3323 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3363 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3682 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3660 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3323 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N490 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4059 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3660 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[11];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6395 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5873 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5846 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5902 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5760, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6434} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5846} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5873} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5902};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6451, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6259} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6395} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5997} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5760};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6388, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6195} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5930} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6305} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6451};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[10];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6015 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6274 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 = !a_man[5];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4053 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3999 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4053 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3631 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3762 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3999 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3631 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3457 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4088 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3415 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3457 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4088 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3839 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3762 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3415 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3954 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3906 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3801 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3954 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3906 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3986 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3242 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4111 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3242 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3833 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3986 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4111 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3962 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3801 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3833 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[8] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3839 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3962 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6532 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[8]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5935, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5744} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6274} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6532};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5931 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6138, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5949} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5935} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6015} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5931};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5987 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5959 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6515, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6327} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5959} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5987} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6056};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5963, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5775} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6138} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6373} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6515};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5897, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6573} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5963} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5820} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6195};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[28], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[27]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6388} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6243} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5897};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7474, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7946} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[28]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[28]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7690, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7676} = {1'B0, N12354} + {1'B0, N12356};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817} = {1'B0, N12294} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7690} + {1'B0, N12298};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3655 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4016 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3655 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4048 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3245 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4016 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4048 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3880 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3977 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3840 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3880 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3977 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3857 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3245 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3840 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4055 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4076 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3597 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4076 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3285 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4055 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3597 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4093 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3474 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4049 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4093 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3474 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3451 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3285 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4049 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N489 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3857 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3451 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6417 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[9];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6502 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6447 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6201, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6011} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6502} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6417} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6447};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6407, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6216} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6201} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5949} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6327};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6333 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6302 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6361 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6310, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6121} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6302} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6333} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6361};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 = !a_man[4];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6331 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 = !a_man[3];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3596 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3217 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3353 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3596 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3217 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3981 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3683 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3945 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3981 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3683 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3431 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3353 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3945 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3547 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3500 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3389 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3547 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3500 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4039 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3582 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4039 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3702 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3423 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3582 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3702 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3553 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3389 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3423 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[6] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3431 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3553 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5778 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[6]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5906, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5723} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6331} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5778};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6069 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[8];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6125 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6001, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5812} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6069} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5906} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6125};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6475 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5871 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3909 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3802 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3909 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3421 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3554 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3802 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3421 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3905 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3252 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3905 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4074 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3882 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4074 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3213 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3252 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3882 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3638 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3554 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3213 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3754 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3704 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3595 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3754 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3704 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3788 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3904 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3632 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3788 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3904 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3761 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3595 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3632 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[7] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3638 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3761 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6151 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[7]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6107, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5921} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5871} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6151};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6392 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5825, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6498} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6107} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6475} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6392};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6087, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5901} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6001} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6121} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6498};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5928 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5898 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5956 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6487, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6295} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5898} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5928} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5956};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5985 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6095 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6012 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6378, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6188} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6095} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5985} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6012};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6579, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6391} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5744} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6487} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6378};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6028, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5840} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6310} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5825} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6434};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5917, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5732} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6579} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6087} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5840};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5852, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6528} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5775} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6407} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5917};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6340, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6148} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5883} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6259} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6028};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[27], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[26]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6340} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5852} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6573};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7548, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7416} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[27]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[27]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7903, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7776} = {1'B0, N12386} + {1'B0, N12388};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420} = {1'B0, N12320} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7903} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7676};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3817 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3844 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3976 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3817 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3844 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3360 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3681 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3360 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3776 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3640 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3681 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3776 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3659 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3976 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3640 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3853 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3390 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4015 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3853 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3390 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3688 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3265 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3845 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3688 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3265 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3244 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4015 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3845 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N488 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3659 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3244 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6037 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6390 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6359 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6414 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6281, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6093} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6359} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6390} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6414};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5888, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6563} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6037} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5921} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6281};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6443 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6556 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6473 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6172, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5984} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6556} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6443} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6473};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6529 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5927 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 = !a_man[2];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 = !a_man[0];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 = !a_man[1];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6387 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6096, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5912} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6387};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6192, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6003} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5927} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6096};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5726 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5798, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6472} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6192} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6529} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5726};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6264, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6076} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5798} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6172} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6295};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6469, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6275} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5888} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6011} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6264};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6499 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[7];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5747 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6549, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6362} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5747} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6499} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5723};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5780, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6454} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6549} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6188} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5812};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5981, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5792} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6391} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5780} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5901};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6292, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6103} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6469} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6216} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5981};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[26], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[25]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6148} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6292} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6528};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7624, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7500} = {1'B0, N12464} + {1'B0, N12466};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7503, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7881} = {1'B0, N12418} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7500};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7624} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7503} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7776};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3400 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3465 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3400 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 = a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3465;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2800 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2820 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2600 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2820} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2800} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2600};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2852 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2830 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2681 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2842 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2704 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2706, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2638} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2842} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2681} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2704};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2830} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2852} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2706};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2771 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2886 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2711 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2747, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2674} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2886} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2771} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2711};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2783 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2783} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2747} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2638};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2745 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2722 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2694 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2649, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2581} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2722} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2745} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2694};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2642 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2630 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2803 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2815 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2878 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2869, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2801} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2815} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2803} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2878};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2791, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2717} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2630} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2642} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2869};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2649} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2674} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2791};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2670 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2790 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2767 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2632, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2883} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2790} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2670} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2767};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2893 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2659 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2734 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2828 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2773, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2699} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2734} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2659} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2828};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2686, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2617} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2893} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2632} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2773};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2581} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2686} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2717};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2593 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2597 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2624 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2713, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2644} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2597} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2593} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2624};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2591, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2843} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2713} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2883} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2699};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2801} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2591} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2617};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2775 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2701 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2811 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2797, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2724} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2701} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2775} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2811};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2781 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2679 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2784 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2666 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2635 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2735, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2665} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2666} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2784} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2635};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2614, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2864} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2679} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2781} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2735};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2671, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2604} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2797} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2644} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2614};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2752 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2844 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2779 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2712 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2602 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2655, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2587} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2712} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2779} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2602};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2853, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2786} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2844} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2752} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2655};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2853} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2671} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2843};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2824 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2838 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2719, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2650} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2824} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2838};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2611 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2708 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2879, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2809} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2611} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2719} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2708};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2753, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2683} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2587} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2724} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2879};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2786} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2753} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2604};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2819 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2850 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2709 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2691 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2805, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2730} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2709} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2691};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2677, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2608} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2850} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2819} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2805};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2647 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2741 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2643 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2858, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2793} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2741} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2647} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2643};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2695, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2623} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2858} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2677} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2665};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2864} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2695} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2683};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2833 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2673 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2829 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2619, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2871} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2673} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2833} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2829};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2826, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2749} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2650} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2619} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2793};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2809} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2826} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2623};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2787 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2877 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2885, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2818} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2787} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2877};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2685 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2891 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2680 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2702, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2633} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2891} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2685} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2680};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2759, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2688} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2885} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2702};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2608} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2759} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2749};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2715 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2732 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2788, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2714} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2715} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2732};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2855 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2845, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2774} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2855} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2788} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2818};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2871} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2845} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2688};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2837 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2867 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2861 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2609 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2595 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2684, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2615} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2609} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2595};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2605, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2854} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2861} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2867} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2684};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2605} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2633} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2774};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2689 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2727 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2578 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2721 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2832, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2754} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2578} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2727} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2721};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2714} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2832} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2854};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2874 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2585 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2778 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2726, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2656} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2585} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2778};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2726} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2615} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2754};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2731 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2616 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2636 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2769, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2616} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2636};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2590 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2590} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2769} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2656};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2682 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2770 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2762 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2629 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2821 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2626, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2629} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2821};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2762} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2770} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2626};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2862 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2723 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2807 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2675 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2807} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2675};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2586 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2763 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2894 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2628 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2763) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2894)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2839 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2868 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2628 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2586) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2839);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2744 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2723) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2868)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2796 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2621 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2744 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2862) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2796);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2846 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2682) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2621)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2661 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2798 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2846 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2731) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2661;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2806 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2576 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2798 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2874) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2806;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2620 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2817 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2576 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2689) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2620;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2761 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2817 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2837) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2761;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2584 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2584;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2720 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2720;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2860 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2860;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2678 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2678;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2827 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2827;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2641 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2641;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2782 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2782;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2599 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2599;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2737 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2737;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2880 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2880;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2696 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2802 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2696;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2588 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174 = N13822 ^ N13824;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[24] = !(N12599 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3341 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3404 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3341 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3436 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3570 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3404 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3436 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3264 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3372 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3226 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3264 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3372 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3243 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3226 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3726 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3447 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3726 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3924 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3614 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3447 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3924 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3272 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3798 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3437 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3272 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3798 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3774 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3614 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3437 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N486 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3243 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3774 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3571 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3259 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3571 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3796 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3796 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3590 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N457 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3259 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3590 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N457;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5152 = !(N14513 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5101 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5217 = !(N12599 | N12753);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5339 = !(N14513 | N12753);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5070 = !(N12599 | N14505);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3751 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3916 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3751 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3371 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3989 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3916 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3371 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3915 = !(a_man[21] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N456 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3989 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3915 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N456;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5272 = !(N13104 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5347, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5270} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5070} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5339} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5272};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[24], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[23]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5217} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5152} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5347};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7523, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7988} = {1'B0, N12538} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[24]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[24]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3615 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3645 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3775 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3615 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3645 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3473 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3572 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3432 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3473 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3572 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3449 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3775 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3432 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3929 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3654 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3929 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4127 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3816 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3654 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4127 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3479 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3995 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3646 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3479 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3995 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3975 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3816 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3646 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N487 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3449 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3975 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6122 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6010 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6181 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6080, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5892} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6010} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6122} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6181};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5954 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4126 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3949 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4083 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4126 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3949 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3780 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3475 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3744 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3780 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3475 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3224 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4083 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3744 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3346 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3487 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3290 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3487 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4125 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3290 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3381 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3498 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3218 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3498 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3352 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4125 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3218 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[5] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3224 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3352 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6262 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5983 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6566, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6382} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6262} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5954} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5983};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6036 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6149 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6065 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6459, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6267} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6149} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6036} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6065};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6061, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5872} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6566} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6080} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6459};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[6];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6233 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6207 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6091 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5971, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5784} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6207} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6233} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6091};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6437, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6247} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6093} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5971} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6472};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6153, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5967} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6061} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6563} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6437};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6495 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5745 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6526 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5877, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6552} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5745} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6495} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6526};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5833 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5806 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6553 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6251, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6064} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5806} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5833} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6553};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5861, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6537} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5877} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6382} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6251};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330 = !(a_man[16] & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3718 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3291 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3543 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3291 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3678 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3718 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3543 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3483 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3377 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3483 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3996 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3336 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3377 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3996 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3756 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3678 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3336 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3871 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3407 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3717 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3871 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3407 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3808 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3907 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3808 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4018 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3747 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3907 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4018 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3876 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3717 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3747 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[3] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3756 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3876 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6376 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[3]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5980 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5920 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6491, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6301} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5980} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6376} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5920};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5724 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5776 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6365, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6177} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5724} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6491} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5776};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6234, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6046} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6365} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5892} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6267};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6329, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6139} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5861} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5872} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6234};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6412 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3923 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3997 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3746 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3997 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3877 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3923 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3746 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4096 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3576 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4096 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3266 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3540 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3576 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3266 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3957 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3877 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3540 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4075 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3619 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3922 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4075 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3619 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4006 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4114 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4006 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3289 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3950 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4114 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3289 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4082 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3922 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3950 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[4] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3957 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4082 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5886 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[4]);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6477, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6284} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5886} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6412} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5912};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6032 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6007 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6063 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6385, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6194} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6007} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6032} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6063};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6178 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[5];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6319 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6230 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5894, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6570} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6319} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6178} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6230};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5767, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6442} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6385} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6284} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5894};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6090 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[4];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6346 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6119 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6270, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6082} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6346} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6090} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6119};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6260 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6204 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6288 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5788, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6461} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6204} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6260} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6288};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6471 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6440 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5858 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5988, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5801} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6440} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6471} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5858};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6143, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5955} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5788} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6270} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5801};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5749, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6425} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5784} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5767} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6143};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6348, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6158} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6477} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6003} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5988};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5952, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5764} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5984} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6348} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6362};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5842, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6517} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6247} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5749} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5764};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6041, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5855} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6329} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5967} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5842};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6534, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6343} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6076} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5952} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6454};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6358, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6167} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6153} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6275} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6534};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[24], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[23]} = {1'B0, N12669} + {1'B0, N12671} + {1'B0, N12673};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[25], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[24]} = {1'B0, N12605} + {1'B0, N12607} + {1'B0, N12609};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7783, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7647} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[24]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[24]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7713, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7972} = {1'B0, N12450} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7523} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7783};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7709, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7568} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[25]} + {1'B0, N12460};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7709} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7713} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7881};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6146 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3517 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3338 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3470 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3338 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3275 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3939 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4110 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3275 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3939 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3799 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4062 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4110 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3799 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3550 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3470 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4062 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3549 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3673 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3549 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3206 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3516 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3673 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3206 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3755 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3705 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3755 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3787 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3819 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3787 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3544 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3705 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3819 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3677 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3516 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3544 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[2] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3550 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3677 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6000 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6436 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6467 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6405, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6213} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6436} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6000} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6467};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6161, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5976} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6405} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6146} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6301};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6521, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6332} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6552} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6161} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6064};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6128, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5938} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6158} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6521} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6537};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5802 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[3];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5970 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5856 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5807, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6481} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5970} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5802} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5856};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6523 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6492 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5914 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5915, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5730} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6492} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6523} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5914};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6551 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5773 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5829 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6290, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6100} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5773} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6551} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5829};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6543, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6352} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5915} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5807} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6290};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5884 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5942 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5743 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6182, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5994} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5942} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5884} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5743};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6051, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5864} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6194} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6182} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6570};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6031, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5845} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6177} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6543} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6051};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6503, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6315} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6046} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6031} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6425};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6218, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6029} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6128} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6139} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6503};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[23], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[22]} = {1'B0, N12744} + {1'B0, N12746} + {1'B0, N12748};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7859, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7730} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[23]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[23]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7922, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7468} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7988} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7647} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7859};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7568} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7922} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7972};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3204 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3804 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3231 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3804 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3370 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3204 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3231 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3270 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3994 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3270 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4104 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3959 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3994 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4104 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3973 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3370 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3959 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3239 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3988 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3719 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3988 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3403 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3239 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3719 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4002 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3592 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3232 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4002 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3592 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3569 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3403 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3232 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N485 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3973 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3569 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5193 = !(N14513 | N14505);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5258 = !(N12599 | N14500);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5125 = !(N13104 | N12753);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5242, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5169} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5258} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5193} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5125};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5316 = !(N13104 | N14505);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5385 = !(N14513 | N14500);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5113 = !(N12599 | N14510);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5330, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5252} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5385} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5316} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5113};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3545 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3575 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3711 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3545 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3575 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3736 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4033 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4103 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4033 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3794 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3711 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4103 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3508 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N455 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3794 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3508 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N455;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5399 = !(N14533 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5390, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5315} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5399} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5330} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5169};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[23], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[22]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5242} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5270} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5390};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7590, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7461} = {1'B0, N12586} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[23]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[23]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3343 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3376 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3509 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3343 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3376 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3534 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3835 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3895 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3534 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3835 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3586 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3509 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3895 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3295 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3868 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3295 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3902 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3301 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3868 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3902 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N454 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3586 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3301 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N454;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5183 = !(N13081 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5247 = !(N14533 | N12753);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5171 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5303 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5235 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5266, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5194} = {1'B0, N13218} + {1'B0, N13220} + {1'B0, N13222};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5141, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5064} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5247} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5183} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5266};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5377 = !(N13081 | N12753);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5104 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4070 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4109 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3302 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4070 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4109 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3327 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3633 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3694 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3327 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3633 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3383 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3302 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3694 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4022 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3668 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4022 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3331 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3700 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3331 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4027 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3668 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3700 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N453 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3383 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4027 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N453;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5308 = !(N14528 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5077, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5341} = {1'B0, N13189} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5377} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5308};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5286, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5211} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5077} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5252} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5064};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[22], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[21]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5141} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5315} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5286};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7940, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7804} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[22]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[22]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7526, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7566} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7461} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7940};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7590} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7526} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7468};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5722 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3274 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3310 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3274 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4066 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3263 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3310 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4066 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4004 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3903 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4004 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3593 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3861 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3903 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3593 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3347 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3263 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3861 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3462 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3940 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3309 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3462 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3940 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3501 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3484 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3581 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3617 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3484 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3581 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3339 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3501 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3617 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3469 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3309 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3339 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[1] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3347 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3469 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6486 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6060 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6086 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6307, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6118} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6060} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6486} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6086};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6557, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6370} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5722} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6213} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6307};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6428, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6240} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6461} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6082} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6557};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6410, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6220} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6442} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6428} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5955};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3411 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4036 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3411 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4124 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3865 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4124 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3992 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3865 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3603 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3701 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3603 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3387 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3662 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3701 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3387 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4079 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3662 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3257 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3739 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4035 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3257 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3739 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3292 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3380 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3405 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3380 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4067 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3292 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3405 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3262 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4035 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4067 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[0] = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4079 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3262 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5841 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6175 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5854 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5828 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5998 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6485, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6294} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5828} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5854} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5998};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6465, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6273} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6175} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5841} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6485};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5960, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5772} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6100} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5994} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6465};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6320, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6131} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6352} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5960} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5864};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5966 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6578 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5881 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5734, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6408} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6578} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5966} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5881};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5741 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[2];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6050 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5913 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6105, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5918} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6050} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5741} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5913};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5979, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5791} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6105} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5734} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6118};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[1];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6079 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5769 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6170 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6199 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6124, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5936} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6170} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6199};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6375, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6186} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5769} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6079} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6124};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5939 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6025 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5800 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5999, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5810} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6025} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5939} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5800};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6374 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6116 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6285 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5822, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6496} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6116} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6374} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6285};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6357, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6165} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5999} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6375} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6496};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6337, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6145} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5979} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6370} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6357};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6144 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6457 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6316 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6197, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6009} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6457} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6144} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6316};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6257 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6227 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6404 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6575, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6389} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6227} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6257} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6404};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6070, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5880} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6575} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6197} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5822};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6344 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6427 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6203 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6084, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5899} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6427} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6344} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6203};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6448, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6256} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6084} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6481};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5944, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5753} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6070} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5976} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6448};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5834, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6509} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6240} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6337} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5753};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6297, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6110} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6320} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5834};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5925, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5736} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6332} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5944} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5845};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6017, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5831} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6410} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5938} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5925};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[21], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[20]} = {1'B0, N12893} + {1'B0, N12895} + {1'B0, N12897};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3733 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3763 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3893 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3733 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3763 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3591 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4030 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3695 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4030 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3551 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3591 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3695 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3567 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3893 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3551 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3770 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3311 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3935 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3770 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3311 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3600 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3461 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3362 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4122 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3461 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3362 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3764 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3600 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4122 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4101 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3935 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3764 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N483 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3567 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4101 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[22], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[21]} = {1'B0, N12823} + {1'B0, N12825} + {1'B0, N12827};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7753, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7612} = {1'B0, N12731} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[21]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[21]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3936 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3964 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4102 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3936 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3964 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3797 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3896 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3758 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3797 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3896 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3773 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4102 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3758 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3970 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3499 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3518 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3499 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3203 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3970 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3518 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3805 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3386 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3965 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3805 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3386 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3369 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3203 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3965 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N484 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3773 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3369 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7673, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7540} = {1'B0, N12647} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[22]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[22]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7734, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7668} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7753} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7804} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7540};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7673} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7734} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7566};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5868, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6545} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6389} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6009} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5899};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5849, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6525} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5880} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5868} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6256};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[0];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6565 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6225 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6254 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5903, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5721} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6225} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6565} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6254};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6513 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6423 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6342 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6500, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6313} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6423} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6513} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6342};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6261, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6073} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6500} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5903} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6294};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6314 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6283 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6371 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6014, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5827} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6283} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6314} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6371};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6516 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6455 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6484 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6399 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6394, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6202} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6484} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6455} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6399};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5885, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6561} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6516} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6014} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6394};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6244, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6055} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5885} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6261} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6273};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6224, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6035} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5772} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6244} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6145};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6209, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6021} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5849} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6131} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6224};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[20], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[19]} = {1'B0, N13000} + {1'B0, N13002} + {1'B0, N13004};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3532 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3555 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3693 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3532 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3555 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4073 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3385 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4073 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3491 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3348 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3385 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3491 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3368 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3693 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3348 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3565 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4019 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4037 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4019 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3732 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3565 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4037 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3391 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3920 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3556 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3391 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3920 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3892 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3732 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3556 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N482 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3368 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3892 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7823, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7698} = {1'B0, N12807} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[20]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[20]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5345 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5279 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5212 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5381, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5305} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5279} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5345} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5212};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3869 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3901 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4028 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3901 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3941 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3424 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3941 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3490 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3424 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4116 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4028 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3490 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3822 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3566 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3458 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3822 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3566 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4057 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3497 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4057 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3830 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3458 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3497 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N452 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4116 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3830 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N452;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5092 = !(N14523 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5353 = !(N14528 | N14505);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5079 = !(N13081 | N14500);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5148 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5187, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5116} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5079} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5353} + {1'B0, N13448};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5356, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5281} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5092} + {1'B0, N13311} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5187};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5087 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5157 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5295 = !(N14533 | N14500);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5398, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5324} = {1'B0, N13335} + {1'B0, N13337} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5295};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3669 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3699 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3831 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3669 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3699 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3652 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3219 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3282 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3652 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3219 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3912 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3831 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3282 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3621 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3365 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3254 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3621 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3365 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3856 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3238 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3288 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3856 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3238 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3629 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3254 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3288 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N451 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3912 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3629 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N451;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5218 = !(N14518 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5284 = !(N14523 | N12753);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5066 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5337 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5215, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5143} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5066} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5337};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5335, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5261} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5284} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5218} + {1'B0, N13424};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5361 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5229 = !(N13081 | N14505);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5162 = !(N14528 | N12753);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5206, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5135} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5229} + {1'B0, N13319} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5162};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5165, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5088} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5335} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5324} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5135};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5374, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5297} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5341} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5356} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5165};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5226, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5153} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5398} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5206} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5194};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[21], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[20]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5226} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5374} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5211};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7408, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7886} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[21]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[21]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7943, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7769} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7823} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7612} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7886};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7408} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7943} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7668};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5777, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6452} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5918} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6408} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5810};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5758, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6433} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5791} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5777} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6165};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6022 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6160 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5922, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5735} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6022} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6160};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6541 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6278, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6089} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6541} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5922} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5936};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6047 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6077 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5995 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6190, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6002} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6077} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6047} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5995};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5910 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5879 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5964 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5814, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6488} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5879} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5910} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5964};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5797 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6104 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5937 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6296, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6109} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6104} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5797} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5937};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5795, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6470} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5814} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6190} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6296};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6150, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5965} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6278} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6186} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5795};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6136 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5824 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5851 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6564, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6380} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5824} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6136} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5851};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6169, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5982} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6564} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5827} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6202};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6530, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6341} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6561} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6169} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6073};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6137, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5948} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6150} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6545} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6530};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5739, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6413} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5758} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6525} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6137};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[19], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[18]} = {1'B0, N13087} + {1'B0, N13089} + {1'B0, N13091};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3326 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3354 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3489 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3326 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3354 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4121 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3283 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4080 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4121 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3283 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4098 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3489 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4080 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3364 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3837 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3531 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3364 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3837 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3585 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4128 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3585 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3716 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3355 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4128 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3716 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3692 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3531 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3355 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N481 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4098 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3692 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7909, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7773} = {1'B0, N12885} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[19]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[19]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5268 = !(N13081 | N14510);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5139 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5071 = !(N14518 | N12753);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5173, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5097} = {1'B0, N13436} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5268} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5071};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5198 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5133 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5204 = !(N14528 | N14500);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5362, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5289} = {1'B0, N13599} + {1'B0, N13601} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5204};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5147, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5073} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5362} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5173} + {1'B0, N13305};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5396 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5260 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3459 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3496 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3630 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3459 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3496 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3444 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3951 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4011 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3444 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3951 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3707 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3630 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4011 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3410 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4095 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3984 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3410 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4095 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3656 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3969 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4017 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3656 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3969 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3419 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3984 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4017 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N450 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3707 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3419 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N450;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5195 = !(N13725 | N12753);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5343, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5267} = {1'B0, N13555} + {1'B0, N13557} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5195};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5122 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5389 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5328 = !(N14523 | N14500);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5196, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5121} = {1'B0, N13591} + {1'B0, N13593} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5328};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5126, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5393} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5196} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5343} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5289};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5312 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5240 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5175 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5223, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5150} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5240} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5312} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5175};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3255 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3287 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3420 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3255 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3287 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3237 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3749 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3813 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3237 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3749 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3505 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3420 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3813 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3209 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3887 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3784 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3209 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3887 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3241 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3768 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3818 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3241 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3768 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3216 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3784 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3818 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N449 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3505 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3216 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N449;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5127 = !(N13712 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5108 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5382 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5245 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5370, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5296} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5382} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5108} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5245};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5155, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5078} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5127} + {1'B0, N13549} + {1'B0, N13551};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5340 = !(N13725 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5254 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5189 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5323 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5387, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5311} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5189} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5254} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5323};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5319, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5244} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5340} + {1'B0, N13430} + {1'B0, N13432};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5273, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5201} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5155} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5097} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5244};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5102, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5368} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5126} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5073} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5273};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5293, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5221} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5319} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5116} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5261};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5310, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5237} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5147} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5281} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5293};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[19], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[18]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5088} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5102} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5237};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[20], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[19]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5153} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5310} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5297};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7561, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7427} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[19]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[19]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7543, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7871} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7909} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7698} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7561};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7489, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7959} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[20]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[20]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7543} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7769};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6482 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5757 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6094, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5909} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6482} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5757};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6367 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6562 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6398 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6474, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6282} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6562} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6367} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6398};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6078, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5889} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6094} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5735} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6474};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6546, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6360} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6313} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5721} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6078};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6453 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6538 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6309 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6363, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6174} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6538} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6453} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6309};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6510 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6339 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6422 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5986, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5799} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6339} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6510} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6422};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6456, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6265} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5986} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6363} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6488};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6058, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5870} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6089} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6456} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6470};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6038, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5853} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6546} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6452} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6058};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6514, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6325} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6055} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6038} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6433};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[18], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[17]} = {1'B0, N13197} + {1'B0, N13199} + {1'B0, N13201};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3782 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4051 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3782 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3402 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4084 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3279 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4051 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4084 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3919 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4012 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3873 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3919 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4012 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3890 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3279 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3873 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4094 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3635 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3325 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4094 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3635 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3925 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3583 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3513 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3583 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4085 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3925 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3513 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3488 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3325 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4085 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N480 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3890 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3488 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7979, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7846} = {1'B0, N12963} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[18]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[18]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7758, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7967} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7979} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7773} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7427};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7959} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7758} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7871};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5733 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6280 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6074 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6217 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5787, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6460} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6074} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6217};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5874, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6550} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6280} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5733} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5787};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5968, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5782} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6109} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6002} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5874};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6435, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6246} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5968} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5982} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6360};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6418, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6228} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5965} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6341} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6435};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[17], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[16]} = {1'B0, N13205} + {1'B0, N13207} + {1'B0, N13209};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3851 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3878 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4008 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3851 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3878 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3715 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3814 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3675 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3715 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3814 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3690 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4008 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3675 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3886 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3426 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4050 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3886 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3426 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3720 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3306 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3879 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3720 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3306 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3278 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4050 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3879 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N479 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3690 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3278 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7450, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7929} = {1'B0, N13074} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[17]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[17]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5386 = !(N13725 | N14505);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5114 = !(N14518 | N14500);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5179 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5177, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5105} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5114} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5386} + {1'B0, N13709};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5318 = !(N13712 | N12753);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5094 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5231 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5395, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5320} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5094} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5231};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5099 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5366 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5299 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5203, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5130} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5366} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5099} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5299};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5326, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5248} = {1'B0, N13689} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5318} + {1'B0, N13693};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5301, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5228} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5177} + {1'B0, N13541} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5326};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5304 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5172 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5220 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5358 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5378, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5302} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5358};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5161, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5084} = {1'B0, N13785} + {1'B0, N13787} + {1'B0, N13789};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5372 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5166 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5236 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5352, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5276} = {1'B0, N13806} + {1'B0, N13808} + {1'B0, N13810};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5137, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5400} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5352} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5161} + {1'B0, N13659};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5111, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5376} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5121} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5267} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5137};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5081, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5349} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5301} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5393} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5111};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[18], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[17]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5221} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5081} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5368};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7637, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7512} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[18]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[18]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7963, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7459} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7450} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7846} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7512};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7637} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7963} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7967};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3650 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3679 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3811 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3650 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3679 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3789 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3512 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3789 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3611 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3466 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3512 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3611 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3485 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3811 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3466 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3972 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3689 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3972 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3222 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3850 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3689 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3222 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3971 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3519 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3971 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4032 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3680 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3519 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4032 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4007 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3850 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3680 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N478 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3485 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4007 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6101 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5933 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6020 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6540, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6350} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5933} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6101} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6020};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5962 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6156 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5992 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6159, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5974} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6156} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5962} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5992};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6249, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6062} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5909} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6540} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6159};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6045 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6132 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6189 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6049, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5862} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6132} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6045} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6189};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5765, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6439} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6049} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5799} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6282};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6345, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6154} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6380} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6249} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5765};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6536 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5813 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5847, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6522} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6536} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5813};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5904 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6426, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6237} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5904} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5847} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6460};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6420 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5754 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6450 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6222, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6034} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5754} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6420} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6450};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6560 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6396 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6479 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5737, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6411} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6396} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6560} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6479};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6507 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5731 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5785 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6113, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5926} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5731} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6507} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5785};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5941, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5751} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5737} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6222} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6113};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6140, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5953} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6174} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6426} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5941};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5857, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6535} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5889} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6265} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6140};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5950, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5762} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6345} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5870} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5857};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[16], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[15]} = {1'B0, N13458} + {1'B0, N13460} + {1'B0, N13462};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7876 = N13094 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[16];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5342 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5145 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5167, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5091} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5342} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5145};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5089 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5144, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5069} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5089} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5167} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5302};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5118, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5384} = {1'B0, N13673} + {1'B0, N13675} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5276};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5090, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5357} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5248} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5118} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5400};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5224 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5154 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5083 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5184, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5112} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5154} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5224} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5083};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5158 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5291 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5363 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5332, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5257} = {1'B0, N13798} + {1'B0, N13800} + {1'B0, N13802};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5307, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5232} = {1'B0, N13697} + {1'B0, N13699} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5332};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5283, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5207} = {1'B0, N13523} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5105} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5307};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5255, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5182} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5078} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5283} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5228};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[16], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[15]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5090} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5376} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5182};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7795, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7663} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[16]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[16]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7564, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7558} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7876} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7929} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7795};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[17], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[16]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5201} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5255} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5349};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7720, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7579} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[17]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[17]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7720} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7564} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7459};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7741 = (!N13094) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[16];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3441 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3471 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3607 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3441 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3471 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3305 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3401 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3260 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3305 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3401 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3276 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3607 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3260 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3481 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3953 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3649 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3481 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3953 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3771 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3312 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3771 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3834 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3472 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3312 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3834 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3810 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3649 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3472 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N477 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3276 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3810 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6318, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6129} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6350} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5974} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5862};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6519, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6330} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6550} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6062} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6318};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6231, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6044} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5782} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6519} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6154};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[15], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[14]} = {1'B0, N13583} + {1'B0, N13585} + {1'B0, N13587};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7602, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7477} = {1'B0, N13466} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[15]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7778, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7662} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7602} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7741} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[16]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7579} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7778} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7558};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5280 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5076 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5214 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5123, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5388} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5076} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5280} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5214};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5346 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5274 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5208 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5313, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5238} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5274} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5346} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5208};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5290, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5216} = {1'B0, N13718} + {1'B0, N13720} + {1'B0, N13722};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5263, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5190} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5084} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5290} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5232};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[15], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[14]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5207} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5263} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5357};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7984, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7762} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7477} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[15]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[15]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7663} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7984} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7662};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6130 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6268 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6287, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6099} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6130} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6268};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6016 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6214 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6040 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5804, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6478} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6214} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6016} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6040};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6490, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6300} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6287} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6522} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5804};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6155 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6187 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6071 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6179, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5991} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6187} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6155} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6071};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6005, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5816} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6179} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6411} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6034};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5832, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6506} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6490} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6237} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6005};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6030, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5844} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6439} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5832} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5953};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[14], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[13]} = {1'B0, N13607} + {1'B0, N13609} + {1'B0, N13611};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6241 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6098 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5728 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5865 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6242, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6053} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5728} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5865};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6555, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6368} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6098} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6241} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6242};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5752 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5811 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6501 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5756, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6431} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5811} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5752} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6501};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6533 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5783 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6558 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6134, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5946} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5783} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6533} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6558};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6067, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5878} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6099} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5756} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6134};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6384, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6193} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6555} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5926} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6067};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6206, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6019} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5751} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6384} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6129};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[13], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[12]} = {1'B0, N13731} + {1'B0, N13733} + {1'B0, N13735};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5067 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5199 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5249 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5391 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5192, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5119} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5249} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5391};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5062, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5327} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5199} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5067} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5192};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5080, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5344} = {1'B0, N13769} + {1'B0, N13771} + {1'B0, N13773};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5129 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5265 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5106, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5371} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5129} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5265};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5134 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5401 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5333 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5250, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5178} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5401} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5134} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5333};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5269, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5197} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5106} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5091} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5250};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5098, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5364} = {1'B0, N13681} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5257} + {1'B0, N13685};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[13], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[12]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5080} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5216} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5364};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7800, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7961} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[13]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[14], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[13]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5098} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5384} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5190};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7585, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7861} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[14]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7456, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7800} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7861};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7456;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7723} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[15]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7585} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7762};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7723;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22792 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6184 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6326 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6572, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6386} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6184} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6326};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5839 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6511, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6322} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5839} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6572} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6053};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6445, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6253} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5991} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6478} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6511};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5893, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6569} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6300} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6445} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5816};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[12], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[11]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6506} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5893} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6019};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5256 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5185 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5120 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5338, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5264} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5256} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5120};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5209, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5138} = {1'B0, N13878} + {1'B0, N13880} + {1'B0, N13882};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[12], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[11]} = {1'B0, N13630} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5209} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5344};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8004, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7452} = {1'B0, N13500} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[12]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8004} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7961};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7997 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6152 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6238 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6293 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6462, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6271} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6238} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6152} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6293};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6211 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6266 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6126 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6083, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5896} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6266} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6211} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6126};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6024, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5837} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6083} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6462} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6431};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5958, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5770} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6368} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6024} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5878};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[11], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[10]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6193} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5958} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6569};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5379 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5176 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5085, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5354} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5379} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5176};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5325 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5151, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5075} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5325} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5085} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5119};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[11], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[10]} = {1'B0, N13761} + {1'B0, N13763} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5138};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7607, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7550} = {1'B0, N13647} + {1'B0, N13649} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[11]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7607} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7452} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[12]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7739 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5809 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5863 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5836 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5929, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5740} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5863} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5809} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5836};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5779 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5919 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6415, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6226} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5779} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5919};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5977, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5789} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6415} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5929} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6386};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6402, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6210} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5946} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5977} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6322};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[10], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[9]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6402} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6253} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5770};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5110 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5309 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5241 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5233, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5309} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5110} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5241};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[10], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[9]} = {1'B0, N13870} + {1'B0, N13872} + {1'B0, N13874};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7819, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7651} = {1'B0, N13777} + {1'B0, N13779} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[10]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7819} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7550};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7476 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5890 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5748 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6232 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6381 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5774, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6449} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6232} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6381};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6304, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6115} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5748} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5890} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5774};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6355, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6162} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5896} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6304} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6271};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[9], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6355} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5837} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6210};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5163 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5300 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5131, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5163} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5300};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5367 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5095 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5287 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5156 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5321, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5287} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5156};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5277, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5095} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5367} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5321};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[9], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5131} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5354} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5277};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7423, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7757} = {1'B0, N13862} + {1'B0, N13864} + {1'B0, N13866};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[10]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7423} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7651};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7814 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6263 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6323 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6291 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6147, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5961} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6323} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6263} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6291};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5819, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6493} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6147} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6226} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5740};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[8], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5819} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5789} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6162};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7631, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7851} = {1'B0, N13896} + {1'B0, N13898} + {1'B0, N13900};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[9]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7631} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7757};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7549 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5916 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5947 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6372, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6183} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5916} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5947};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6351 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6527, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6338} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6351} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6372} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6449};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[7], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6527} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6115} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6493};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7839, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7949} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[7]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974} = {1'B0, N13835} + {1'B0, N13837} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7851};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7902 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5859 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5887 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5975 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5882, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5887} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5859} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5975};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[6], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[5]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5882} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5961} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6338};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[6] = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7445, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7444} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[6]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574} = {1'B0, N13888} + {1'B0, N13890} + {1'B0, N13892};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7625 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[5] = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6377 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6406 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6483, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[3]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6377} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6406};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6430 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6347 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5969 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6027 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6102, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[2]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5969} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6027};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5996, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[3]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6347} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6430} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6102};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[5], float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6483} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6183} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5996};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[5] = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7656, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7546} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[5]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7925, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7789} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7656} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7444};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7969 = !(N13842 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[4] = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7868, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7642} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[4]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[4]};
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7528, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7868} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7546};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7711 = N13854 & N13856;
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[4]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7642};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7436 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[3]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[3]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7786 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[2] = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531);
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547, float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7414} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[2]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[2]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7525 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7895 = !(((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7636 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7895 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7414);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7990 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7487 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7636 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7525) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7990);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7857 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7786) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7487)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7921 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7623 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7857 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7436) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7921);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7926 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7711) & (!N13852)) | ((!N13854) & (!N13856));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7831 = !(N13842 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7609 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7926 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7969) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7831);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7828 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7625) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7609)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7763 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7442 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7828 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7902) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7763);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7583 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7549) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7442)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7688 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7733 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7583 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7814) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7688);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7796 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7476) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7733)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7599 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7860 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7796 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7739) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7599);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7694 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7997) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7860)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7552 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22792) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7694)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11605 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11605 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7552) | (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005) | (!(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934) | (!(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853) | (!(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779) | (!(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703) | (!(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620) | (!(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544) | (!(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593)) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467 = N12206 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467) | (!(N12206 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415)) | ((!N12194) & (!N12196));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7993 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7692 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854 & N11929) | (!(N12176 | N12178)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438 = ((!N12097) & (!N12095)) | ((!N12184) & (!N12186));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7924 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775 ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438 & N12092) | (!(N12166 | N12168)));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486 = ((!N12087) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806)) | ((!N12144) & (!N12146));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486 | (!N12082));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7970 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768 | N12077) & (N12110 | N12112);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7889 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3894 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7790 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3894 | a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7765 = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7889) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7790;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[39] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7970) ^ N12072;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2523 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2514 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2526 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2518 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2516 = !(((float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2523 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2514) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2526) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2518);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2516 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[7] = !a_exp[7];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[5] = !a_exp[5];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[3] = !a_exp[3];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[1] = !a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[0] = !a_exp[0];
assign {float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[0]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[0]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0]};
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[1] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457 = !(a_exp[2] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[3] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451 = !(a_exp[4] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[5] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444 = !(a_exp[6] & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[2] = (!a_exp[2]) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[3] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[3]) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[5] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[5]) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2486 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[2] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[3]) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[6] = (!a_exp[6]) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[7] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[7]) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2489 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[6] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[4] = (!a_exp[4]) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[1] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[1]) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2483 = !((((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2489) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[0]) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[4]) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N446 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2486 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2483);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__17 = ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444) & (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[7])) | (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N446);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N447 = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__17);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33 = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29 | (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N447));
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_N448 = ((float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0] | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__67 = !float_div_cynw_cm_float_rcp_E8_M23_2_inst_N448;
assign x[22] = (N12012 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[39]) | ((!N12012) & N12014);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[38] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768) ^ N12077;
assign x[21] = (N12012 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[38]) | ((!N12012) & N12014);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[37] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486) ^ N12082;
assign x[20] = (N12012 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[37]) | ((!N12012) & N12014);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[36] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806) ^ N12087;
assign x[19] = (N12012 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[36]) | ((!N12012) & N12014);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[35] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438) ^ N12092;
assign x[18] = (N12012 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[35]) | ((!N12012) & N12014);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[34] = (!N12095) ^ N12097;
assign x[17] = (N12012 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[34]) | ((!N12012) & N12014);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[33] = (!N13225) ^ N13227;
assign x[16] = (N12012 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[33]) | ((!N12012) & N12014);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[32] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[15] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[32]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[31] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[14] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[31]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[30] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[13] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[30]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[29] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[12] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[29]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[28] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[11] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[28]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[27] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[10] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[27]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[26] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[9] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[26]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[25] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[8] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[25]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[24] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[7] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[24]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[23] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[6] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[23]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[22] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[5] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[22]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[21] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[4] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[21]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[20] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[3] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[20]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[19] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[2] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[19]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[18] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[1] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[18]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[17] = (!float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002) ^ float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[0] = (N11736 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[17]) | ((!N11736) & N11738);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38 = float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 = !((float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34) | float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[30] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[7]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[29] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[6]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[28] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[5]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[27] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[4]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[26] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[3]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[25] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[2]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[24] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[1]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[23] = (float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[0]) | ((!float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[31] = !(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29 | (!a_sign));
reg x_reg_L0_23__I2241_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__I2241_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[23];
	end
assign N5603 = x_reg_L0_23__I2241_QOUT;
reg x_reg_L0_24__I2242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_24__I2242_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[24];
	end
assign N5608 = x_reg_L0_24__I2242_QOUT;
reg x_reg_L0_25__I2243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_25__I2243_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[25];
	end
assign N5613 = x_reg_L0_25__I2243_QOUT;
reg x_reg_L0_26__I2244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_26__I2244_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[26];
	end
assign N5618 = x_reg_L0_26__I2244_QOUT;
reg x_reg_L0_27__I2245_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_27__I2245_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[27];
	end
assign N5623 = x_reg_L0_27__I2245_QOUT;
reg x_reg_L0_28__I2246_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_28__I2246_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[28];
	end
assign N5628 = x_reg_L0_28__I2246_QOUT;
reg x_reg_L0_29__I2247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_29__I2247_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[29];
	end
assign N5633 = x_reg_L0_29__I2247_QOUT;
reg x_reg_L0_30__I2248_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_30__I2248_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[30];
	end
assign N5638 = x_reg_L0_30__I2248_QOUT;
reg x_reg_L0_31__I2249_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__I2249_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[31];
	end
assign N5643 = x_reg_L0_31__I2249_QOUT;
reg x_reg_L1_0__I2250_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__I2250_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[0];
	end
assign x[0] = x_reg_L1_0__I2250_QOUT;
reg x_reg_L1_1__I2251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__I2251_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[1];
	end
assign x[1] = x_reg_L1_1__I2251_QOUT;
reg x_reg_L1_2__I2252_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__I2252_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[2];
	end
assign x[2] = x_reg_L1_2__I2252_QOUT;
reg x_reg_L1_3__I2253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__I2253_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[3];
	end
assign x[3] = x_reg_L1_3__I2253_QOUT;
reg x_reg_L1_4__I2254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__I2254_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[4];
	end
assign x[4] = x_reg_L1_4__I2254_QOUT;
reg x_reg_L1_5__I2255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__I2255_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[5];
	end
assign x[5] = x_reg_L1_5__I2255_QOUT;
reg x_reg_L1_6__I2256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__I2256_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[6];
	end
assign x[6] = x_reg_L1_6__I2256_QOUT;
reg x_reg_L1_7__I2257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__I2257_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[7];
	end
assign x[7] = x_reg_L1_7__I2257_QOUT;
reg x_reg_L1_8__I2258_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__I2258_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[8];
	end
assign x[8] = x_reg_L1_8__I2258_QOUT;
reg x_reg_L1_9__I2259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__I2259_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[9];
	end
assign x[9] = x_reg_L1_9__I2259_QOUT;
reg x_reg_L1_10__I2260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__I2260_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[10];
	end
assign x[10] = x_reg_L1_10__I2260_QOUT;
reg x_reg_L1_11__I2261_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__I2261_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[11];
	end
assign x[11] = x_reg_L1_11__I2261_QOUT;
reg x_reg_L1_12__I2262_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__I2262_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[12];
	end
assign x[12] = x_reg_L1_12__I2262_QOUT;
reg x_reg_L1_13__I2263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__I2263_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[13];
	end
assign x[13] = x_reg_L1_13__I2263_QOUT;
reg x_reg_L1_14__I2264_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__I2264_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[14];
	end
assign x[14] = x_reg_L1_14__I2264_QOUT;
reg x_reg_L1_15__I2265_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__I2265_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[15];
	end
assign x[15] = x_reg_L1_15__I2265_QOUT;
reg x_reg_L1_23__I2273_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__I2273_QOUT <= N5603;
	end
assign x[23] = x_reg_L1_23__I2273_QOUT;
reg x_reg_L1_24__I2274_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__I2274_QOUT <= N5608;
	end
assign x[24] = x_reg_L1_24__I2274_QOUT;
reg x_reg_L1_25__I2275_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__I2275_QOUT <= N5613;
	end
assign x[25] = x_reg_L1_25__I2275_QOUT;
reg x_reg_L1_26__I2276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__I2276_QOUT <= N5618;
	end
assign x[26] = x_reg_L1_26__I2276_QOUT;
reg x_reg_L1_27__I2277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__I2277_QOUT <= N5623;
	end
assign x[27] = x_reg_L1_27__I2277_QOUT;
reg x_reg_L1_28__I2278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__I2278_QOUT <= N5628;
	end
assign x[28] = x_reg_L1_28__I2278_QOUT;
reg x_reg_L1_29__I2279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__I2279_QOUT <= N5633;
	end
assign x[29] = x_reg_L1_29__I2279_QOUT;
reg x_reg_L1_30__I2280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__I2280_QOUT <= N5638;
	end
assign x[30] = x_reg_L1_30__I2280_QOUT;
reg x_reg_L1_31__I2281_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I2281_QOUT <= N5643;
	end
assign x[31] = x_reg_L1_31__I2281_QOUT;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[16] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  vLfwTgnbqhs= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



