/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:25:15 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_3 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__9,
	inst_cellmath__10,
	inst_cellmath__11,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__16,
	inst_cellmath__17,
	inst_cellmath__18;
wire [8:0] inst_cellmath__27,
	inst_cellmath__28;
wire [7:0] inst_cellmath__29;
wire  inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__32;
wire [49:0] inst_cellmath__33;
wire  inst_cellmath__34;
wire [7:0] inst_cellmath__35;
wire [49:0] inst_cellmath__36,
	inst_cellmath__37;
wire [25:0] inst_cellmath__39;
wire  inst_cellmath__42,
	inst_cellmath__43,
	inst_cellmath__44;
wire [26:0] inst_cellmath__45;
wire  inst_cellmath__48;
wire [5:0] inst_cellmath__49;
wire [24:0] inst_cellmath__50;
wire  inst_cellmath__53,
	inst_cellmath__54,
	inst_cellmath__55;
wire [23:0] inst_cellmath__57;
wire [9:0] inst_cellmath__59;
wire  inst_cellmath__62,
	inst_cellmath__63;
wire [22:0] inst_cellmath__64;
wire  inst_cellmath__66;
wire [7:0] inst_cellmath__68;
wire  inst_cellmath__70;
wire N547,N556,N557,N558,N559,N560,N561 
	,N562,N563,N565,N567,N568,N569,N570,N571 
	,N572,N574,N575,N625,N626,N627,N628,N630 
	,N631,N632,N633,N634,N635,N636,N638,N639 
	,N642,N645,N650,N651,N652,N653,N655,N656 
	,N657,N658,N659,N660,N661,N662,N663,N664 
	,N665,N666,N667,N668,N669,N670,N671,N672 
	,N673,N674,N675,N676,N677,N706,N710,N2691 
	,N4132,N4134,N4155,N4163,N4166,N4168,N4172,N4174 
	,N4177,N4183,N4187,N4218,N4221,N4232,N4240,N4243 
	,N4245,N4249,N4251,N4254,N4260,N4264,N4310,N4314 
	,N4336,N4340,N4357,N4360,N4364,N4368,N4370,N4372 
	,N4373,N4375,N4376,N4377,N4379,N4380,N4382,N4384 
	,N4386,N4387,N4390,N4393,N4396,N4401,N4402,N4404 
	,N4405,N4407,N4408,N4414,N4417,N4418,N4466,N4467 
	,N4468,N4469,N4471,N4473,N4475,N4476,N4477,N4478 
	,N4479,N4482,N4483,N4484,N4486,N4487,N4489,N4491 
	,N4493,N4494,N4495,N4496,N4497,N4499,N4500,N4502 
	,N4504,N4506,N4507,N4509,N4510,N4512,N4514,N4516 
	,N4517,N4518,N4520,N4522,N4523,N4524,N4525,N4528 
	,N4530,N4531,N4533,N4534,N4536,N4538,N4540,N4541 
	,N4542,N4543,N4545,N4546,N4548,N4550,N4551,N4552 
	,N4553,N4555,N4557,N4558,N4559,N4561,N4562,N4564 
	,N4565,N4566,N4567,N4568,N4569,N4570,N4571,N4574 
	,N4575,N4576,N4578,N4580,N4581,N4583,N4585,N4587 
	,N4588,N4590,N4591,N4593,N4595,N4597,N4598,N4599 
	,N4600,N4602,N4603,N4604,N4605,N4607,N4609,N4610 
	,N4611,N4613,N4614,N4751,N4792,N4793,N4832,N4903 
	,N4905,N4906,N4907,N4909,N4911,N4912,N4914,N4915 
	,N4916,N4918,N4920,N4921,N4922,N4923,N4925,N4927 
	,N4929,N4930,N4931,N4932,N4935,N4937,N4939,N4940 
	,N4942,N4944,N4946,N4947,N4948,N4949,N4952,N4953 
	,N4954,N4955,N4956,N4958,N4959,N4960,N4962,N4964 
	,N4965,N4967,N4969,N4970,N4972,N4974,N4976,N4977 
	,N4978,N4979,N4982,N4983,N4984,N4986,N4988,N4989 
	,N4990,N4991,N4993,N4995,N4997,N4998,N5000,N5002 
	,N5003,N5005,N5008,N5010,N5012,N5013,N5014,N5015 
	,N5017,N5019,N5021,N5022,N5023,N5025,N5027,N5028 
	,N5029,N5031,N5033,N5034,N5036,N5038,N5040,N5041 
	,N5042,N5043,N5046,N5047,N5048,N5049,N5051,N5053 
	,N5055,N5056,N5057,N5059,N5061,N5062,N5064,N5066 
	,N5068,N5069,N5070,N5071,N5074,N5075,N5077,N5079 
	,N5080,N5081,N5082,N5084,N5085,N5087,N5089,N5090 
	,N5092,N5094,N5095,N5096,N5097,N5098,N5100,N5103 
	,N5104,N5105,N5107,N5109,N5110,N5111,N5112,N5114 
	,N5116,N5119,N5120,N5342,N5397,N5398,N5400,N5402 
	,N5404,N5407,N5408,N5411,N5414,N5416,N5418,N5419 
	,N5421,N5427,N5428,N5431,N5436,N5437,N5465,N5643 
	,N5644,N5646,N5648,N5650,N5651,N5652,N5655,N5656 
	,N5657,N5659,N5660,N5661,N5664,N5665,N5666,N5667 
	,N5668,N5671,N5672,N5674,N5675,N5677,N5679,N5680 
	,N5682,N5684,N5686,N5687,N5689,N5691,N5693,N5694 
	,N5695,N5698,N5700,N5701,N5702,N5703,N5706,N5707 
	,N5708,N5710,N5711,N5714,N5715,N5717,N5718,N5721 
	,N5723,N5724,N5725,N5728,N5730,N5731,N5734,N5735 
	,N5737,N5738,N5741,N5742,N5744,N5745,N5746,N5749 
	,N5750,N5752,N5753,N5756,N5758,N5759,N5760,N5763 
	,N5765,N5766,N5767,N5770,N5771,N5772,N5773,N5775 
	,N5777,N5778,N5779,N5781,N5783,N5785,N5786,N5788 
	,N5790,N5791,N5792,N5793,N5796,N5798,N5800,N5801 
	,N5803,N5805,N5806,N5808,N5809,N5811,N5813,N5814 
	,N5816,N5817,N5819,N5820,N5822,N5823,N5824,N5827 
	,N5829,N5830,N5831,N5832,N5835,N5836,N5837,N5838 
	,N5839,N5840,N5993,N5995,N5996,N5997,N5998,N6000 
	,N6001,N6004,N6005,N6006,N6007,N6009,N6010,N6011 
	,N6014,N6015,N6016,N6017,N6019,N6021,N6024,N6025 
	,N6026,N6028,N6029,N6031,N6032,N6033,N6035,N6037 
	,N6038,N6039,N6041,N6042,N6043,N6046,N6047,N6049 
	,N6050,N6052,N6054,N6056,N6057,N6058,N6060,N6061 
	,N6062,N6063,N6065,N6067,N6069,N6070,N6071,N6073 
	,N6074,N6076,N6078,N6079,N6080,N6082,N6083,N6086 
	,N6087,N6212,N6233,N6282,N6285,N6291,N6297,N6298 
	,N6300,N6301,N6303,N6306,N6307,N6308,N6310,N6311 
	,N6312,N6314,N6315,N6317,N6318,N6319,N6321,N6323 
	,N6324,N6326,N6328,N6330,N6331,N6333,N6334,N6335 
	,N6337,N6338,N6341,N6343,N6344,N6346,N6347,N6349 
	,N6350,N6352,N6353,N6355,N6357,N6358,N6360,N6361 
	,N6362,N6364,N6365,N6367,N6368,N6371,N6373,N6374 
	,N6375,N6377,N6379,N6380,N6382,N6383,N6385,N6386 
	,N6387,N6389,N6390,N6392,N6394,N6395,N6397,N6398 
	,N6400,N6402,N6404,N6405,N6407,N6408,N6409,N6411 
	,N6412,N6414,N6416,N6417,N6419,N6420,N6422,N6423 
	,N6424,N6426,N6427,N6429,N6430,N6432,N6434,N6435 
	,N6436,N6438,N6439,N6441,N6443,N6444,N6445,N6447 
	,N6448,N6450,N6452,N6453,N6454,N6456,N6457,N6459 
	,N6460,N6655,N6695,N6696,N6701,N6702,N6703,N6705 
	,N6709,N6710,N6713,N6714,N6718,N6719,N6720,N6721 
	,N6727,N6729,N6731,N6732,N6734,N6744,N6748,N6749 
	,N6751,N6754,N6758,N6759,N6762,N6763,N6766,N6767 
	,N6768,N6769,N6770,N6775,N6776,N6777,N6883,N6889 
	,N6892,N6893,N6901,N6902,N6905,N6908,N6909,N6911 
	,N6913,N6917,N6918,N6919,N6921,N6923,N6928,N6929 
	,N6930,N6931,N6932,N6933,N6936,N6938,N6941,N6944 
	,N6946,N6948,N6950,N6951,N6954,N6997,N6999,N7000 
	,N7018,N7020,N7056,N7068,N7074,N7092,N7111,N7117 
	,N7122,N7125,N7129,N7133,N7138,N7141,N7142,N7146 
	,N7150,N7153,N7156,N7161,N7166,N7169,N7173,N7178 
	,N7182,N7186,N7190,N7195,N7198,N7202,N7207,N7210 
	,N8708,N8722,N8730,N8733,N8738,N8749,N8772,N8785 
	,N8801,N8804,N8806,N8808,N8809,N8812,N8814,N8816 
	,N8817,N8820,N8824,N8825,N8826,N8830,N8834,N8840 
	,N8847,N8854,N8861,N8868,N8875,N8882,N13892,N13893 
	,N13895;
XOR2XL cynw_cm_float_add2_ieee_I706 (.Y(inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
NAND2XL inst_cellmath__9_0_I707 (.Y(N4132), .A(a_exp[0]), .B(a_exp[1]));
AND4XL inst_cellmath__9_0_I7910 (.Y(N4134), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3282 (.Y(N8834), .A(a_exp[7]), .B(a_exp[6]), .C(N4134));
NOR2XL hyperpropagate_4_1_A_I3283 (.Y(inst_cellmath__9), .A(N4132), .B(N8834));
NOR2XL inst_cellmath__10__1__I720 (.Y(N4155), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__10__1__I721 (.Y(N4163), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__10__1__I722 (.Y(N4174), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__10__1__I723 (.Y(N4183), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__10__1__I7911 (.Y(N4168), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__10__1__I7912 (.Y(N4177), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__10__1__I7913 (.Y(N4187), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__10__1__I727 (.Y(N4172), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N4168));
NAND4XL inst_cellmath__10__1__I729 (.Y(N4166), .A(N4155), .B(N4174), .C(N4163), .D(N4183));
NOR4BX1 inst_cellmath__10__1__I7914 (.Y(inst_cellmath__10), .AN(N4172), .B(N4166), .C(N4177), .D(N4187));
AND2XL cynw_cm_float_add2_ieee_I732 (.Y(inst_cellmath__12), .A(inst_cellmath__9), .B(inst_cellmath__10));
NAND4XL inst_cellmath__14_0_I733 (.Y(N4221), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[7]), .D(b_exp[6]));
INVXL cynw_cm_float_add2_ieee_I18 (.Y(N559), .A(b_exp[3]));
INVXL cynw_cm_float_add2_ieee_I424 (.Y(N2691), .A(N559));
NAND4XL inst_cellmath__14_0_I734 (.Y(N4218), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[2]), .D(N2691));
NOR2XL inst_cellmath__14_0_I735 (.Y(inst_cellmath__14), .A(N4221), .B(N4218));
NOR2XL inst_cellmath__15__3__I742 (.Y(N4232), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__15__3__I743 (.Y(N4240), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__15__3__I744 (.Y(N4251), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__15__3__I745 (.Y(N4260), .A(b_man[4]), .B(b_man[3]));
OR4X1 inst_cellmath__15__3__I7915 (.Y(N4245), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__15__3__I7916 (.Y(N4254), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__15__3__I7917 (.Y(N4264), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4X1 inst_cellmath__15__3__I749 (.Y(N4249), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N4245));
NAND4XL inst_cellmath__15__3__I751 (.Y(N4243), .A(N4232), .B(N4251), .C(N4240), .D(N4260));
NOR4BX1 inst_cellmath__15__3__I7918 (.Y(inst_cellmath__15), .AN(N4249), .B(N4243), .C(N4254), .D(N4264));
AND2XL cynw_cm_float_add2_ieee_I754 (.Y(inst_cellmath__17), .A(inst_cellmath__15), .B(inst_cellmath__14));
AND3XL cynw_cm_float_add2_ieee_I755 (.Y(N547), .A(inst_cellmath__12), .B(inst_cellmath__17), .C(inst_cellmath__39[25]));
NOR2BX1 cynw_cm_float_add2_ieee_I756 (.Y(inst_cellmath__13), .AN(inst_cellmath__9), .B(inst_cellmath__10));
NOR2BX1 cynw_cm_float_add2_ieee_I757 (.Y(inst_cellmath__18), .AN(inst_cellmath__14), .B(inst_cellmath__15));
OR3XL cynw_cm_float_add2_ieee_I758 (.Y(inst_cellmath__63), .A(inst_cellmath__13), .B(inst_cellmath__18), .C(N547));
OR4X1 inst_cellmath__11__2__I7919 (.Y(N4310), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 inst_cellmath__11__2__I7920 (.Y(N4314), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL inst_cellmath__11__2__I765 (.Y(inst_cellmath__11), .A(N4310), .B(N4314));
OR4X1 inst_cellmath__16__4__I7921 (.Y(N4340), .A(b_exp[7]), .B(b_exp[5]), .C(b_exp[6]), .D(b_exp[4]));
OR4X1 inst_cellmath__16__4__I769 (.Y(N4336), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[2]), .D(N2691));
NOR2XL inst_cellmath__16__4__I770 (.Y(inst_cellmath__16), .A(N4340), .B(N4336));
AND2XL cynw_cm_float_add2_ieee_I771 (.Y(N706), .A(inst_cellmath__11), .B(inst_cellmath__16));
NOR3BXL cynw_cm_float_add2_ieee_I772 (.Y(inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
INVXL cynw_cm_float_add2_ieee_I15 (.Y(N556), .A(b_exp[0]));
INVX2 cynw_cm_float_add2_ieee_I16 (.Y(N557), .A(b_exp[1]));
INVXL cynw_cm_float_add2_ieee_I17 (.Y(N558), .A(b_exp[2]));
INVXL cynw_cm_float_add2_ieee_I19 (.Y(N560), .A(b_exp[4]));
INVXL cynw_cm_float_add2_ieee_I20 (.Y(N561), .A(b_exp[5]));
INVXL cynw_cm_float_add2_ieee_I21 (.Y(N562), .A(b_exp[6]));
INVXL cynw_cm_float_add2_ieee_I22 (.Y(N563), .A(b_exp[7]));
NAND2XL inst_cellmath__28__8__I773 (.Y(N4404), .A(a_exp[0]), .B(N556));
OR2XL inst_cellmath__28__8__I774 (.Y(N4372), .A(a_exp[1]), .B(N557));
INVX1 inst_cellmath__28__8__I3074 (.Y(N8733), .A(a_exp[1]));
MXI2X1 inst_cellmath__28__8__I3075 (.Y(N8730), .A(a_exp[1]), .B(N8733), .S0(N557));
INVX1 inst_cellmath__28__8__I3076 (.Y(N4364), .A(N8730));
NOR2XL inst_cellmath__28__8__I776 (.Y(N4380), .A(a_exp[2]), .B(N558));
XOR2XL inst_cellmath__28__8__I777 (.Y(N4396), .A(a_exp[2]), .B(N558));
OR2XL inst_cellmath__28__8__I778 (.Y(N4377), .A(a_exp[3]), .B(N559));
XOR2XL inst_cellmath__28__8__I779 (.Y(N4360), .A(a_exp[3]), .B(N559));
OR2XL inst_cellmath__28__8__I780 (.Y(N4417), .A(a_exp[4]), .B(N560));
XOR2XL inst_cellmath__28__8__I781 (.Y(N4386), .A(a_exp[4]), .B(N560));
OR2XL inst_cellmath__28__8__I782 (.Y(N4382), .A(a_exp[5]), .B(N561));
XOR2XL inst_cellmath__28__8__I783 (.Y(N4418), .A(a_exp[5]), .B(N561));
OR2XL inst_cellmath__28__8__I784 (.Y(N4357), .A(a_exp[6]), .B(N562));
XOR2XL inst_cellmath__28__8__I785 (.Y(N4376), .A(a_exp[6]), .B(N562));
NOR2XL inst_cellmath__28__8__I786 (.Y(N4393), .A(a_exp[7]), .B(N563));
XOR2XL inst_cellmath__28__8__I787 (.Y(N4408), .A(a_exp[7]), .B(N563));
OAI2BB1X1 inst_cellmath__28__8__I788 (.Y(N4384), .A0N(N4364), .A1N(N4404), .B0(N4372));
INVXL gen2_alt_A_I3284 (.Y(N8840), .A(N4380));
OAI2BB1X1 gen2_alt_A_I3285 (.Y(N4405), .A0N(N4396), .A1N(N4384), .B0(N8840));
OAI2BB1XL inst_cellmath__28__8__I791 (.Y(N4387), .A0N(N4360), .A1N(N4405), .B0(N4377));
OAI2BB1XL inst_cellmath__28__8__I792 (.Y(N4401), .A0N(N4386), .A1N(N4387), .B0(N4417));
OAI2BB1XL inst_cellmath__28__8__I793 (.Y(N4370), .A0N(N4418), .A1N(N4401), .B0(N4382));
OAI2BB1XL inst_cellmath__28__8__I794 (.Y(N4375), .A0N(N4376), .A1N(N4370), .B0(N4357));
XOR2XL inst_cellmath__28__8__I796 (.Y(N565), .A(a_exp[0]), .B(N556));
XNOR2X1 inst_cellmath__28__8__I3077 (.Y(N8738), .A(N4404), .B(N4364));
XNOR2X1 inst_cellmath__28__8__I798 (.Y(N567), .A(N4384), .B(N4396));
XNOR2X1 inst_cellmath__28__8__I799 (.Y(N568), .A(N4405), .B(N4360));
XNOR2X1 inst_cellmath__28__8__I800 (.Y(N569), .A(N4387), .B(N4386));
XNOR2X1 inst_cellmath__28__8__I801 (.Y(N570), .A(N4401), .B(N4418));
XNOR2X1 inst_cellmath__28__8__I802 (.Y(N571), .A(N4370), .B(N4376));
XNOR2X1 inst_cellmath__28__8__I803 (.Y(N572), .A(N4375), .B(N4408));
NOR2XL inst_cellmath__28__8__I804 (.Y(N4368), .A(N556), .B(a_exp[0]));
OAI2BB1X1 inst_cellmath__28__8__I805 (.Y(N4407), .A0N(N4368), .A1N(N4364), .B0(N4372));
INVXL gen2_alt_A_I3286 (.Y(N8847), .A(N4380));
OAI2BB1X1 gen2_alt_A_I3287 (.Y(N4390), .A0N(N4396), .A1N(N4407), .B0(N8847));
OAI2BB1XL inst_cellmath__28__8__I807 (.Y(N4402), .A0N(N4360), .A1N(N4390), .B0(N4377));
OAI2BB1XL inst_cellmath__28__8__I808 (.Y(N4373), .A0N(N4386), .A1N(N4402), .B0(N4417));
OAI2BB1XL inst_cellmath__28__8__I809 (.Y(N4379), .A0N(N4418), .A1N(N4373), .B0(N4382));
OAI2BB1X1 inst_cellmath__28__8__I810 (.Y(N4414), .A0N(N4376), .A1N(N4379), .B0(N4357));
INVXL gen2_alt_A_I3288 (.Y(N8854), .A(N4393));
OAI2BB1X1 gen2_alt_A_I3289 (.Y(inst_cellmath__27[8]), .A0N(N4408), .A1N(N4414), .B0(N8854));
BUFX3 inst_cellmath__28__8__I3200 (.Y(N8801), .A(inst_cellmath__27[8]));
XOR2XL inst_cellmath__28__8__I812 (.Y(inst_cellmath__27[0]), .A(a_exp[0]), .B(N556));
XOR2XL inst_cellmath__28__8__I813 (.Y(inst_cellmath__27[1]), .A(N4368), .B(N4364));
XOR2XL inst_cellmath__28__8__I814 (.Y(inst_cellmath__27[2]), .A(N4407), .B(N4396));
XOR2XL inst_cellmath__28__8__I815 (.Y(inst_cellmath__27[3]), .A(N4390), .B(N4360));
XOR2XL inst_cellmath__28__8__I816 (.Y(inst_cellmath__27[4]), .A(N4402), .B(N4386));
XOR2XL inst_cellmath__28__8__I817 (.Y(inst_cellmath__27[5]), .A(N4373), .B(N4418));
XOR2XL inst_cellmath__28__8__I818 (.Y(inst_cellmath__27[6]), .A(N4379), .B(N4376));
XOR2XL inst_cellmath__28__8__I819 (.Y(inst_cellmath__27[7]), .A(N4414), .B(N4408));
AOI21X1 cynw_cm_float_add2_ieee_I3100 (.Y(inst_cellmath__28[8]), .A0(N4408), .A1(N4375), .B0(N4393));
INVXL inst_cellmath__34_0_I820 (.Y(N4497), .A(a_man[1]));
INVXL inst_cellmath__34_0_I821 (.Y(N4564), .A(a_man[2]));
INVXL inst_cellmath__34_0_I822 (.Y(N4478), .A(a_man[3]));
INVXL inst_cellmath__34_0_I823 (.Y(N4543), .A(a_man[4]));
INVXL inst_cellmath__34_0_I824 (.Y(N4610), .A(a_man[5]));
INVXL inst_cellmath__34_0_I825 (.Y(N4524), .A(a_man[6]));
INVXL inst_cellmath__34_0_I826 (.Y(N4588), .A(a_man[7]));
INVXL inst_cellmath__34_0_I827 (.Y(N4507), .A(a_man[8]));
INVXL inst_cellmath__34_0_I828 (.Y(N4570), .A(a_man[9]));
INVXL inst_cellmath__34_0_I829 (.Y(N4484), .A(a_man[10]));
INVXL inst_cellmath__34_0_I830 (.Y(N4552), .A(a_man[11]));
INVXL inst_cellmath__34_0_I831 (.Y(N4468), .A(a_man[12]));
INVXL inst_cellmath__34_0_I832 (.Y(N4531), .A(a_man[13]));
INVXL inst_cellmath__34_0_I833 (.Y(N4598), .A(a_man[14]));
INVXL inst_cellmath__34_0_I834 (.Y(N4516), .A(a_man[15]));
INVXL inst_cellmath__34_0_I835 (.Y(N4578), .A(a_man[16]));
INVXL inst_cellmath__34_0_I836 (.Y(N4494), .A(a_man[17]));
INVXL inst_cellmath__34_0_I837 (.Y(N4561), .A(a_man[18]));
INVXL inst_cellmath__34_0_I838 (.Y(N4473), .A(a_man[19]));
INVXL inst_cellmath__34_0_I839 (.Y(N4541), .A(a_man[20]));
INVXL inst_cellmath__34_0_I840 (.Y(N4607), .A(a_man[21]));
INVXL inst_cellmath__34_0_I841 (.Y(N4520), .A(a_man[22]));
INVXL inst_cellmath__34_0_I842 (.Y(N4504), .A(b_man[0]));
NAND2XL inst_cellmath__34_0_I843 (.Y(N4512), .A(b_man[1]), .B(N4497));
NOR2XL inst_cellmath__34_0_I844 (.Y(N4477), .A(b_man[1]), .B(N4497));
NAND2XL inst_cellmath__34_0_I845 (.Y(N4609), .A(b_man[2]), .B(N4564));
NOR2XL inst_cellmath__34_0_I846 (.Y(N4575), .A(b_man[2]), .B(N4564));
NAND2XL inst_cellmath__34_0_I847 (.Y(N4557), .A(b_man[3]), .B(N4478));
NOR2XL inst_cellmath__34_0_I848 (.Y(N4523), .A(b_man[3]), .B(N4478));
NAND2XL inst_cellmath__34_0_I849 (.Y(N4506), .A(b_man[4]), .B(N4543));
NOR2XL inst_cellmath__34_0_I850 (.Y(N4471), .A(b_man[4]), .B(N4543));
NAND2XL inst_cellmath__34_0_I851 (.Y(N4603), .A(b_man[5]), .B(N4610));
NOR2XL inst_cellmath__34_0_I852 (.Y(N4569), .A(b_man[5]), .B(N4610));
NAND2XL inst_cellmath__34_0_I853 (.Y(N4551), .A(b_man[6]), .B(N4524));
NOR2XL inst_cellmath__34_0_I854 (.Y(N4518), .A(b_man[6]), .B(N4524));
NAND2XL inst_cellmath__34_0_I855 (.Y(N4500), .A(b_man[7]), .B(N4588));
NOR2XL inst_cellmath__34_0_I856 (.Y(N4467), .A(b_man[7]), .B(N4588));
NAND2XL inst_cellmath__34_0_I857 (.Y(N4597), .A(b_man[8]), .B(N4507));
NOR2XL inst_cellmath__34_0_I858 (.Y(N4566), .A(b_man[8]), .B(N4507));
NAND2XL inst_cellmath__34_0_I859 (.Y(N4546), .A(b_man[9]), .B(N4570));
NOR2XL inst_cellmath__34_0_I860 (.Y(N4514), .A(b_man[9]), .B(N4570));
NAND2XL inst_cellmath__34_0_I861 (.Y(N4493), .A(b_man[10]), .B(N4484));
NOR2XL inst_cellmath__34_0_I862 (.Y(N4613), .A(b_man[10]), .B(N4484));
NAND2XL inst_cellmath__34_0_I863 (.Y(N4591), .A(b_man[11]), .B(N4552));
NOR2XL inst_cellmath__34_0_I864 (.Y(N4559), .A(b_man[11]), .B(N4552));
NAND2XL inst_cellmath__34_0_I865 (.Y(N4540), .A(b_man[12]), .B(N4468));
NOR2XL inst_cellmath__34_0_I866 (.Y(N4509), .A(b_man[12]), .B(N4468));
NAND2XL inst_cellmath__34_0_I867 (.Y(N4487), .A(b_man[13]), .B(N4531));
NOR2XL inst_cellmath__34_0_I868 (.Y(N4605), .A(b_man[13]), .B(N4531));
NAND2XL inst_cellmath__34_0_I869 (.Y(N4587), .A(b_man[14]), .B(N4598));
NOR2XL inst_cellmath__34_0_I870 (.Y(N4555), .A(b_man[14]), .B(N4598));
NAND2XL inst_cellmath__34_0_I871 (.Y(N4534), .A(b_man[15]), .B(N4516));
NOR2XL inst_cellmath__34_0_I872 (.Y(N4502), .A(b_man[15]), .B(N4516));
NAND2XL inst_cellmath__34_0_I873 (.Y(N4482), .A(b_man[16]), .B(N4578));
NOR2XL inst_cellmath__34_0_I874 (.Y(N4600), .A(b_man[16]), .B(N4578));
NAND2XL inst_cellmath__34_0_I875 (.Y(N4581), .A(b_man[17]), .B(N4494));
NOR2XL inst_cellmath__34_0_I876 (.Y(N4548), .A(b_man[17]), .B(N4494));
NAND2XL inst_cellmath__34_0_I877 (.Y(N4528), .A(b_man[18]), .B(N4561));
NOR2XL inst_cellmath__34_0_I878 (.Y(N4496), .A(b_man[18]), .B(N4561));
NAND2XL inst_cellmath__34_0_I879 (.Y(N4476), .A(b_man[19]), .B(N4473));
NOR2XL inst_cellmath__34_0_I880 (.Y(N4593), .A(b_man[19]), .B(N4473));
NAND2XL inst_cellmath__34_0_I881 (.Y(N4574), .A(b_man[20]), .B(N4541));
NOR2XL inst_cellmath__34_0_I882 (.Y(N4542), .A(b_man[20]), .B(N4541));
NAND2XL inst_cellmath__34_0_I883 (.Y(N4522), .A(b_man[21]), .B(N4607));
NOR2XL inst_cellmath__34_0_I884 (.Y(N4489), .A(b_man[21]), .B(N4607));
OR2XL inst_cellmath__34_0_I885 (.Y(N4538), .A(b_man[22]), .B(N4520));
OAI21XL inst_cellmath__34_0_I886 (.Y(N4536), .A0(N4489), .A1(N4574), .B0(N4522));
NOR2XL inst_cellmath__34_0_I887 (.Y(N4568), .A(N4489), .B(N4542));
OAI21XL inst_cellmath__34_0_I888 (.Y(N4602), .A0(N4593), .A1(N4528), .B0(N4476));
NOR2XL inst_cellmath__34_0_I889 (.Y(N4483), .A(N4593), .B(N4496));
OAI21XL inst_cellmath__34_0_I890 (.Y(N4517), .A0(N4548), .A1(N4482), .B0(N4581));
NOR2XL inst_cellmath__34_0_I891 (.Y(N4550), .A(N4548), .B(N4600));
OAI21XL inst_cellmath__34_0_I892 (.Y(N4583), .A0(N4502), .A1(N4587), .B0(N4534));
NOR2XL inst_cellmath__34_0_I893 (.Y(N4466), .A(N4502), .B(N4555));
OAI21XL inst_cellmath__34_0_I894 (.Y(N4499), .A0(N4605), .A1(N4540), .B0(N4487));
NOR2XL inst_cellmath__34_0_I895 (.Y(N4530), .A(N4605), .B(N4509));
OAI21XL inst_cellmath__34_0_I896 (.Y(N4565), .A0(N4559), .A1(N4493), .B0(N4591));
NOR2XL inst_cellmath__34_0_I897 (.Y(N4595), .A(N4559), .B(N4613));
OAI21XL inst_cellmath__34_0_I898 (.Y(N4479), .A0(N4514), .A1(N4597), .B0(N4546));
OAI21XL inst_cellmath__34_0_I900 (.Y(N4545), .A0(N4467), .A1(N4551), .B0(N4500));
NOR2XL inst_cellmath__34_0_I901 (.Y(N4576), .A(N4467), .B(N4518));
OAI21XL inst_cellmath__34_0_I902 (.Y(N4611), .A0(N4569), .A1(N4506), .B0(N4603));
NOR2XL inst_cellmath__34_0_I903 (.Y(N4491), .A(N4569), .B(N4471));
OAI21XL inst_cellmath__34_0_I904 (.Y(N4525), .A0(N4523), .A1(N4609), .B0(N4557));
NOR2XL inst_cellmath__34_0_I905 (.Y(N4558), .A(N4523), .B(N4575));
OAI31X1 inst_cellmath__34_0_I906 (.Y(N4590), .A0(N4504), .A1(a_man[0]), .A2(N4477), .B0(N4512));
AOI22XL inst_cellmath__34_0_I907 (.Y(N4571), .A0(N4538), .A1(N4536), .B0(b_man[22]), .B1(N4520));
NAND2XL inst_cellmath__34_0_I908 (.Y(N4604), .A(N4538), .B(N4568));
AOI21XL inst_cellmath__34_0_I909 (.Y(N4486), .A0(N4483), .A1(N4517), .B0(N4602));
AOI21XL inst_cellmath__34_0_I910 (.Y(N4553), .A0(N4466), .A1(N4499), .B0(N4583));
NAND2XL inst_cellmath__34_0_I911 (.Y(N4585), .A(N4466), .B(N4530));
AOI21XL inst_cellmath__34_0_I912 (.Y(N4469), .A0(N4595), .A1(N4479), .B0(N4565));
NOR4BX1 inst_cellmath__34_0_I7925 (.Y(N4614), .AN(N4595), .B(N4514), .C(N4585), .D(N4566));
AOI21XL inst_cellmath__34_0_I914 (.Y(N4533), .A0(N4576), .A1(N4611), .B0(N4545));
NAND2XL inst_cellmath__34_0_I915 (.Y(N4567), .A(N4576), .B(N4491));
AOI21XL inst_cellmath__34_0_I916 (.Y(N4599), .A0(N4558), .A1(N4590), .B0(N4525));
NAND3BXL inst_cellmath__34_0_I917 (.Y(N4510), .AN(N4604), .B(N4483), .C(N4550));
OAI21XL inst_cellmath__34_0_I918 (.Y(N4580), .A0(N4585), .A1(N4469), .B0(N4553));
OAI21XL inst_cellmath__34_0_I920 (.Y(N4495), .A0(N4567), .A1(N4599), .B0(N4533));
AOI21XL inst_cellmath__34_0_I921 (.Y(N4562), .A0(N4614), .A1(N4495), .B0(N4580));
OA21X1 inst_cellmath__34_0_I922 (.Y(N4475), .A0(N4604), .A1(N4486), .B0(N4571));
OAI21XL inst_cellmath__34_0_I923 (.Y(inst_cellmath__34), .A0(N4510), .A1(N4562), .B0(N4475));
NOR2BX1 cynw_cm_float_add2_ieee_I924 (.Y(N575), .AN(inst_cellmath__34), .B(inst_cellmath__28[8]));
NOR2X1 cynw_cm_float_add2_ieee_I925 (.Y(inst_cellmath__32), .A(inst_cellmath__27[8]), .B(N575));
MX2XL cynw_cm_float_add2_ieee_I926 (.Y(inst_cellmath__48), .A(b_sign), .B(a_sign), .S0(inst_cellmath__32));
INVX3 inst_cellmath__35_0_I935 (.Y(N4751), .A(N8801));
AOI22X2 inst_cellmath__35_0_I936 (.Y(inst_cellmath__35[0]), .A0(N4751), .A1(inst_cellmath__27[0]), .B0(N565), .B1(N8801));
AOI22X2 inst_cellmath__35_0_I3080 (.Y(N8749), .A0(inst_cellmath__27[1]), .A1(N4751), .B0(N8738), .B1(N8801));
AOI22X1 inst_cellmath__35_0_I938 (.Y(inst_cellmath__35[2]), .A0(inst_cellmath__27[2]), .A1(N4751), .B0(N567), .B1(N8801));
AOI22XL inst_cellmath__35_0_I939 (.Y(inst_cellmath__35[3]), .A0(N4751), .A1(inst_cellmath__27[3]), .B0(N568), .B1(N8801));
AOI22XL inst_cellmath__35_0_I940 (.Y(inst_cellmath__35[4]), .A0(N4751), .A1(inst_cellmath__27[4]), .B0(N569), .B1(N8801));
AOI22XL inst_cellmath__35_0_I941 (.Y(inst_cellmath__35[5]), .A0(N4751), .A1(inst_cellmath__27[5]), .B0(N570), .B1(N8801));
AOI22XL inst_cellmath__35_0_I942 (.Y(inst_cellmath__35[6]), .A0(N4751), .A1(inst_cellmath__27[6]), .B0(N571), .B1(N8801));
AOI22XL inst_cellmath__35_0_I943 (.Y(inst_cellmath__35[7]), .A0(N4751), .A1(inst_cellmath__27[7]), .B0(N572), .B1(N8801));
OAI211X1 inst_cellmath__30_0_I944 (.Y(N4793), .A0(inst_cellmath__35[2]), .A1(N8749), .B0(inst_cellmath__35[4]), .C0(inst_cellmath__35[3]));
NOR3BXL inst_cellmath__30_0_I945 (.Y(N4792), .AN(N4793), .B(inst_cellmath__35[6]), .C(inst_cellmath__35[5]));
NAND2BXL inst_cellmath__30_0_I946 (.Y(inst_cellmath__30), .AN(inst_cellmath__35[7]), .B(N4792));
OR2XL cynw_cm_float_add2_ieee_I947 (.Y(inst_cellmath__31), .A(inst_cellmath__11), .B(inst_cellmath__16));
CLKINVX6 inst_cellmath__36__15__I950 (.Y(N4832), .A(inst_cellmath__32));
MX2XL inst_cellmath__36__15__I951 (.Y(inst_cellmath__36[26]), .A(b_man[0]), .B(a_man[0]), .S0(N4832));
MX2XL inst_cellmath__36__15__I952 (.Y(inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(N4832));
MX2XL inst_cellmath__36__15__I953 (.Y(inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(N4832));
MX2XL inst_cellmath__36__15__I954 (.Y(inst_cellmath__36[29]), .A(b_man[3]), .B(a_man[3]), .S0(N4832));
MX2XL inst_cellmath__36__15__I955 (.Y(inst_cellmath__36[30]), .A(b_man[4]), .B(a_man[4]), .S0(N4832));
MX2XL inst_cellmath__36__15__I956 (.Y(inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(N4832));
MX2XL inst_cellmath__36__15__I957 (.Y(inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(N4832));
MX2XL inst_cellmath__36__15__I958 (.Y(inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(N4832));
MX2XL inst_cellmath__36__15__I959 (.Y(inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(N4832));
MX2XL inst_cellmath__36__15__I960 (.Y(inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(N4832));
MX2XL inst_cellmath__36__15__I961 (.Y(inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(N4832));
MX2XL inst_cellmath__36__15__I962 (.Y(inst_cellmath__36[37]), .A(b_man[11]), .B(a_man[11]), .S0(N4832));
MX2XL inst_cellmath__36__15__I963 (.Y(inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(N4832));
MX2XL inst_cellmath__36__15__I964 (.Y(inst_cellmath__36[39]), .A(b_man[13]), .B(a_man[13]), .S0(N4832));
MX2XL inst_cellmath__36__15__I965 (.Y(inst_cellmath__36[40]), .A(b_man[14]), .B(a_man[14]), .S0(N4832));
MX2XL inst_cellmath__36__15__I966 (.Y(inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(N4832));
MX2XL inst_cellmath__36__15__I967 (.Y(inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(N4832));
MX2XL inst_cellmath__36__15__I3201 (.Y(inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(N4832));
MX2XL inst_cellmath__36__15__I969 (.Y(inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(N4832));
MX2XL inst_cellmath__36__15__I970 (.Y(inst_cellmath__36[45]), .A(b_man[19]), .B(a_man[19]), .S0(N4832));
MX2XL inst_cellmath__36__15__I971 (.Y(inst_cellmath__36[46]), .A(b_man[20]), .B(a_man[20]), .S0(N4832));
MX2XL inst_cellmath__36__15__I972 (.Y(inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(N4832));
MX2XL inst_cellmath__36__15__I973 (.Y(inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(N4832));
INVX3 inst_cellmath__37_0_I974 (.Y(N5084), .A(inst_cellmath__35[0]));
NOR2BX1 inst_cellmath__37_0_I975 (.Y(N4955), .AN(inst_cellmath__36[26]), .B(N5084));
MX2XL inst_cellmath__37_0_I976 (.Y(N5048), .A(inst_cellmath__36[27]), .B(inst_cellmath__36[26]), .S0(N5084));
MX2XL inst_cellmath__37_0_I977 (.Y(N5096), .A(inst_cellmath__36[28]), .B(inst_cellmath__36[27]), .S0(N5084));
MX2XL inst_cellmath__37_0_I978 (.Y(N4930), .A(inst_cellmath__36[29]), .B(inst_cellmath__36[28]), .S0(N5084));
MX2XL inst_cellmath__37_0_I979 (.Y(N4978), .A(inst_cellmath__36[30]), .B(inst_cellmath__36[29]), .S0(N5084));
MX2XL inst_cellmath__37_0_I980 (.Y(N5022), .A(inst_cellmath__36[31]), .B(inst_cellmath__36[30]), .S0(N5084));
MX2XL inst_cellmath__37_0_I981 (.Y(N5069), .A(inst_cellmath__36[32]), .B(inst_cellmath__36[31]), .S0(N5084));
MX2XL inst_cellmath__37_0_I982 (.Y(N5120), .A(inst_cellmath__36[33]), .B(inst_cellmath__36[32]), .S0(N5084));
MX2XL inst_cellmath__37_0_I983 (.Y(N4947), .A(inst_cellmath__36[34]), .B(inst_cellmath__36[33]), .S0(N5084));
MX2XL inst_cellmath__37_0_I984 (.Y(N4998), .A(inst_cellmath__36[35]), .B(inst_cellmath__36[34]), .S0(N5084));
MX2XL inst_cellmath__37_0_I985 (.Y(N5042), .A(inst_cellmath__36[36]), .B(inst_cellmath__36[35]), .S0(N5084));
MX2XL inst_cellmath__37_0_I986 (.Y(N5090), .A(inst_cellmath__36[37]), .B(inst_cellmath__36[36]), .S0(N5084));
MX2XL inst_cellmath__37_0_I987 (.Y(N4921), .A(inst_cellmath__36[38]), .B(inst_cellmath__36[37]), .S0(N5084));
MX2XL inst_cellmath__37_0_I988 (.Y(N4970), .A(inst_cellmath__36[39]), .B(inst_cellmath__36[38]), .S0(N5084));
MX2XL inst_cellmath__37_0_I989 (.Y(N5013), .A(inst_cellmath__36[40]), .B(inst_cellmath__36[39]), .S0(N5084));
MX2XL inst_cellmath__37_0_I990 (.Y(N5062), .A(inst_cellmath__36[41]), .B(inst_cellmath__36[40]), .S0(N5084));
MX2XL inst_cellmath__37_0_I991 (.Y(N5110), .A(inst_cellmath__36[42]), .B(inst_cellmath__36[41]), .S0(N5084));
MX2XL inst_cellmath__37_0_I992 (.Y(N4940), .A(inst_cellmath__36[43]), .B(inst_cellmath__36[42]), .S0(N5084));
MX2XL inst_cellmath__37_0_I993 (.Y(N4989), .A(inst_cellmath__36[44]), .B(inst_cellmath__36[43]), .S0(N5084));
MX2XL inst_cellmath__37_0_I994 (.Y(N5034), .A(inst_cellmath__36[45]), .B(inst_cellmath__36[44]), .S0(N5084));
MX2XL inst_cellmath__37_0_I995 (.Y(N5080), .A(inst_cellmath__36[46]), .B(inst_cellmath__36[45]), .S0(N5084));
MX2XL inst_cellmath__37_0_I996 (.Y(N4912), .A(inst_cellmath__36[47]), .B(inst_cellmath__36[46]), .S0(N5084));
MX2XL inst_cellmath__37_0_I997 (.Y(N4959), .A(inst_cellmath__36[48]), .B(inst_cellmath__36[47]), .S0(N5084));
NAND2BXL inst_cellmath__37_0_I998 (.Y(N5005), .AN(inst_cellmath__36[48]), .B(N5084));
INVX2 inst_cellmath__37_0_I999 (.Y(N4914), .A(inst_cellmath__35[2]));
INVX2 inst_cellmath__37_0_I1000 (.Y(N4964), .A(N4914));
NAND2XL inst_cellmath__37_0_I1001 (.Y(N5103), .A(N4964), .B(N4955));
NAND2XL inst_cellmath__37_0_I1002 (.Y(N4982), .A(N4964), .B(N5048));
NAND2XL inst_cellmath__37_0_I1003 (.Y(N5074), .A(N4964), .B(N5096));
NAND2XL inst_cellmath__37_0_I1004 (.Y(N4952), .A(N4964), .B(N4930));
AOI22XL inst_cellmath__37_0_I1005 (.Y(N5046), .A0(N4964), .A1(N4978), .B0(N4955), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1006 (.Y(N5094), .A0(N4964), .A1(N5022), .B0(N5048), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1007 (.Y(N4927), .A0(N4964), .A1(N5069), .B0(N5096), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1008 (.Y(N4974), .A0(N4964), .A1(N5120), .B0(N4930), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1009 (.Y(N5019), .A0(N4964), .A1(N4947), .B0(N4978), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1010 (.Y(N5066), .A0(N4964), .A1(N4998), .B0(N5022), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1011 (.Y(N5116), .A0(N4964), .A1(N5042), .B0(N5069), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1012 (.Y(N4944), .A0(N4964), .A1(N5090), .B0(N5120), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1013 (.Y(N4995), .A0(N4964), .A1(N4921), .B0(N4947), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1014 (.Y(N5038), .A0(N4964), .A1(N4970), .B0(N4998), .B1(N4914));
AOI22X1 inst_cellmath__37_0_I1015 (.Y(N5087), .A0(N4964), .A1(N5013), .B0(N5042), .B1(N4914));
AOI22XL inst_cellmath__37_0_I3137 (.Y(N4918), .A0(N4914), .A1(N5090), .B0(N4964), .B1(N5062));
AOI22XL inst_cellmath__37_0_I1017 (.Y(N4967), .A0(N4964), .A1(N5110), .B0(N4921), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1018 (.Y(N5010), .A0(N4964), .A1(N4940), .B0(N4970), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1019 (.Y(N5059), .A0(N4964), .A1(N4989), .B0(N5013), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1020 (.Y(N5107), .A0(N4964), .A1(N5034), .B0(N5062), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1021 (.Y(N4937), .A0(N4964), .A1(N5080), .B0(N5110), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1022 (.Y(N4986), .A0(N4964), .A1(N4912), .B0(N4940), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1023 (.Y(N5031), .A0(N4964), .A1(N4959), .B0(N4989), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1024 (.Y(N5077), .A0(N4964), .A1(N5005), .B0(N5034), .B1(N4914));
AOI22XL inst_cellmath__37_0_I1025 (.Y(N4909), .A0(N5084), .A1(N4964), .B0(N5080), .B1(N4914));
NAND2XL inst_cellmath__37_0_I1026 (.Y(N4956), .A(N4912), .B(N4914));
NAND2XL inst_cellmath__37_0_I1027 (.Y(N5049), .A(N4959), .B(N4914));
NAND2XL inst_cellmath__37_0_I1028 (.Y(N4931), .A(N5005), .B(N4914));
NAND2XL inst_cellmath__37_0_I1029 (.Y(N5023), .A(N5084), .B(N4914));
INVX1 inst_cellmath__37_0_I1030 (.Y(N5055), .A(N8749));
INVX1 inst_cellmath__37_0_I1031 (.Y(N5104), .A(N5055));
NOR2XL inst_cellmath__37_0_I1032 (.Y(N4915), .A(N5055), .B(N5103));
NOR2XL inst_cellmath__37_0_I1033 (.Y(N5056), .A(N5055), .B(N4982));
AOI22XL inst_cellmath__37_0_I1034 (.Y(N4984), .A0(N5055), .A1(N5103), .B0(N5074), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1035 (.Y(N5028), .A0(N5055), .A1(N4982), .B0(N4952), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1036 (.Y(N5075), .A0(N5055), .A1(N5074), .B0(N5046), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1037 (.Y(N4906), .A0(N5055), .A1(N4952), .B0(N5094), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1038 (.Y(N4954), .A0(N5055), .A1(N5046), .B0(N4927), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1039 (.Y(N5002), .A0(N5055), .A1(N5094), .B0(N4974), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1040 (.Y(N5047), .A0(N5055), .A1(N4927), .B0(N5019), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1041 (.Y(N5095), .A0(N5055), .A1(N4974), .B0(N5066), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1042 (.Y(N4929), .A0(N5055), .A1(N5019), .B0(N5116), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1043 (.Y(N4976), .A0(N5055), .A1(N5066), .B0(N4944), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1044 (.Y(N5021), .A0(N5055), .A1(N5116), .B0(N4995), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1045 (.Y(N5068), .A0(N5055), .A1(N4944), .B0(N5038), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1046 (.Y(N5119), .A0(N5055), .A1(N4995), .B0(N5087), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1047 (.Y(N4946), .A0(N5055), .A1(N5038), .B0(N4918), .B1(N5104));
AOI22X1 inst_cellmath__37_0_I1048 (.Y(N4997), .A0(N5055), .A1(N5087), .B0(N4967), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1049 (.Y(N5040), .A0(N5055), .A1(N4918), .B0(N5010), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1050 (.Y(N5089), .A0(N5055), .A1(N4967), .B0(N5059), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1051 (.Y(N4920), .A0(N5055), .A1(N5010), .B0(N5107), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1052 (.Y(N4969), .A0(N5055), .A1(N5059), .B0(N4937), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1053 (.Y(N5012), .A0(N5055), .A1(N5107), .B0(N4986), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1054 (.Y(N5061), .A0(N5055), .A1(N4937), .B0(N5031), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1055 (.Y(N5109), .A0(N5055), .A1(N4986), .B0(N5077), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1056 (.Y(N4939), .A0(N5055), .A1(N5031), .B0(N4909), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1057 (.Y(N4988), .A0(N5055), .A1(N5077), .B0(N4956), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1058 (.Y(N5033), .A0(N5055), .A1(N4909), .B0(N5049), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1059 (.Y(N5079), .A0(N5055), .A1(N4956), .B0(N4931), .B1(N5104));
AOI22XL inst_cellmath__37_0_I1060 (.Y(N4911), .A0(N5055), .A1(N5049), .B0(N5023), .B1(N5104));
NOR2XL inst_cellmath__37_0_I1061 (.Y(N4958), .A(N5104), .B(N4931));
NOR2XL inst_cellmath__37_0_I1062 (.Y(N5100), .A(N5104), .B(N5023));
INVX1 inst_cellmath__37_0_I1063 (.Y(N4983), .A(inst_cellmath__35[4]));
INVX1 inst_cellmath__37_0_I1064 (.Y(N5027), .A(N4983));
NAND2XL inst_cellmath__37_0_I1065 (.Y(N5098), .A(N5027), .B(N4915));
NAND2XL inst_cellmath__37_0_I1066 (.Y(N4979), .A(N5027), .B(N5056));
NAND2XL inst_cellmath__37_0_I1067 (.Y(N5071), .A(N5027), .B(N4984));
NAND2XL inst_cellmath__37_0_I1068 (.Y(N4949), .A(N5027), .B(N5028));
NAND2XL inst_cellmath__37_0_I1069 (.Y(N5043), .A(N5027), .B(N5075));
NAND2XL inst_cellmath__37_0_I1070 (.Y(N4923), .A(N5027), .B(N4906));
NAND2XL inst_cellmath__37_0_I1071 (.Y(N5015), .A(N5027), .B(N4954));
NAND2XL inst_cellmath__37_0_I1072 (.Y(N5112), .A(N5027), .B(N5002));
NAND2XL inst_cellmath__37_0_I1073 (.Y(N4991), .A(N5027), .B(N5047));
NAND2XL inst_cellmath__37_0_I1074 (.Y(N5082), .A(N5027), .B(N5095));
NAND2XL inst_cellmath__37_0_I1075 (.Y(N4962), .A(N5027), .B(N4929));
NAND2XL inst_cellmath__37_0_I1076 (.Y(N5053), .A(N5027), .B(N4976));
NAND2XL inst_cellmath__37_0_I1077 (.Y(N4932), .A(N5027), .B(N5021));
NAND2XL inst_cellmath__37_0_I1078 (.Y(N5025), .A(N5027), .B(N5068));
NAND2XL inst_cellmath__37_0_I1079 (.Y(N4903), .A(N5027), .B(N5119));
NAND2XL inst_cellmath__37_0_I1080 (.Y(N5000), .A(N5027), .B(N4946));
AOI22XL inst_cellmath__37_0_I1081 (.Y(N5092), .A0(N5027), .A1(N4997), .B0(N4915), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1082 (.Y(N4925), .A0(N5027), .A1(N5040), .B0(N5056), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1083 (.Y(N4972), .A0(N5027), .A1(N5089), .B0(N4984), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1084 (.Y(N5017), .A0(N5027), .A1(N4920), .B0(N5028), .B1(N4983));
AOI22XL inst_cellmath__37_0_I3105 (.Y(N5064), .A0(N4983), .A1(N5075), .B0(N5027), .B1(N4969));
AOI22XL inst_cellmath__37_0_I1086 (.Y(N5114), .A0(N5027), .A1(N5012), .B0(N4906), .B1(N4983));
AOI22XL inst_cellmath__37_0_I3106 (.Y(N4942), .A0(N4983), .A1(N4954), .B0(N5027), .B1(N5061));
AOI22XL inst_cellmath__37_0_I1088 (.Y(N4993), .A0(N5027), .A1(N5109), .B0(N5002), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1089 (.Y(N5036), .A0(N5027), .A1(N4939), .B0(N5047), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1090 (.Y(N5085), .A0(N5027), .A1(N4988), .B0(N5095), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1091 (.Y(N4916), .A0(N5027), .A1(N5033), .B0(N4929), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1092 (.Y(N4965), .A0(N5027), .A1(N5079), .B0(N4976), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1093 (.Y(N5008), .A0(N5027), .A1(N4911), .B0(N5021), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1094 (.Y(N5057), .A0(N5027), .A1(N4958), .B0(N5068), .B1(N4983));
AOI22XL inst_cellmath__37_0_I1095 (.Y(N5105), .A0(N5027), .A1(N5100), .B0(N5119), .B1(N4983));
NAND2XL inst_cellmath__37_0_I1096 (.Y(N4935), .A(N4946), .B(N4983));
NAND2XL inst_cellmath__37_0_I1097 (.Y(N5029), .A(N4997), .B(N4983));
NAND2XL inst_cellmath__37_0_I1098 (.Y(N4907), .A(N5040), .B(N4983));
NAND2XL inst_cellmath__37_0_I1099 (.Y(N5003), .A(N5089), .B(N4983));
NAND2XL inst_cellmath__37_0_I3203 (.Y(N5097), .A(N4920), .B(N4983));
NAND2XL inst_cellmath__37_0_I1101 (.Y(N4977), .A(N4969), .B(N4983));
NAND2XL inst_cellmath__37_0_I1102 (.Y(N5070), .A(N5012), .B(N4983));
NAND2XL inst_cellmath__37_0_I1103 (.Y(N4948), .A(N5061), .B(N4983));
NAND2XL inst_cellmath__37_0_I1104 (.Y(N5041), .A(N5109), .B(N4983));
NAND2XL inst_cellmath__37_0_I1105 (.Y(N4922), .A(N4939), .B(N4983));
NAND2XL inst_cellmath__37_0_I1106 (.Y(N5014), .A(N4988), .B(N4983));
NAND2XL inst_cellmath__37_0_I1107 (.Y(N5111), .A(N5033), .B(N4983));
NAND2XL inst_cellmath__37_0_I1108 (.Y(N4990), .A(N5079), .B(N4983));
NAND2XL inst_cellmath__37_0_I1109 (.Y(N5081), .A(N4911), .B(N4983));
NAND2XL inst_cellmath__37_0_I1110 (.Y(N4960), .A(N4958), .B(N4983));
NAND2XL inst_cellmath__37_0_I1111 (.Y(N5051), .A(N5100), .B(N4983));
INVX2 inst_cellmath__37_0_I3204 (.Y(N4905), .A(inst_cellmath__35[3]));
INVX1 inst_cellmath__37_0_I1114 (.Y(N4953), .A(N4905));
NOR2XL inst_cellmath__37_0_I1115 (.Y(inst_cellmath__37[0]), .A(N4905), .B(N4923));
NOR2X1 inst_cellmath__37_0_I1116 (.Y(inst_cellmath__37[1]), .A(N4905), .B(N5015));
NOR2XL inst_cellmath__37_0_I1117 (.Y(inst_cellmath__37[2]), .A(N4905), .B(N5112));
AOI22XL inst_cellmath__37_0_I1118 (.Y(inst_cellmath__37[3]), .A0(N4905), .A1(N5098), .B0(N4991), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1119 (.Y(inst_cellmath__37[4]), .A0(N4905), .A1(N4979), .B0(N5082), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1120 (.Y(inst_cellmath__37[5]), .A0(N4905), .A1(N5071), .B0(N4962), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1121 (.Y(inst_cellmath__37[6]), .A0(N4905), .A1(N4949), .B0(N5053), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1122 (.Y(inst_cellmath__37[7]), .A0(N4905), .A1(N5043), .B0(N4932), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1123 (.Y(inst_cellmath__37[8]), .A0(N4905), .A1(N4923), .B0(N5025), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1124 (.Y(inst_cellmath__37[9]), .A0(N4905), .A1(N5015), .B0(N4903), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1125 (.Y(inst_cellmath__37[10]), .A0(N4905), .A1(N5112), .B0(N5000), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1126 (.Y(inst_cellmath__37[11]), .A0(N4905), .A1(N4991), .B0(N5092), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1127 (.Y(inst_cellmath__37[12]), .A0(N4905), .A1(N5082), .B0(N4925), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1128 (.Y(inst_cellmath__37[13]), .A0(N4905), .A1(N4962), .B0(N4972), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1129 (.Y(inst_cellmath__37[14]), .A0(N4905), .A1(N5053), .B0(N5017), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1130 (.Y(inst_cellmath__37[15]), .A0(N4905), .A1(N4932), .B0(N5064), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1131 (.Y(inst_cellmath__37[16]), .A0(N4905), .A1(N5025), .B0(N5114), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1132 (.Y(inst_cellmath__37[17]), .A0(N4905), .A1(N4903), .B0(N4942), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1133 (.Y(inst_cellmath__37[18]), .A0(N4905), .A1(N5000), .B0(N4993), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1134 (.Y(inst_cellmath__37[19]), .A0(N4905), .A1(N5092), .B0(N5036), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1135 (.Y(inst_cellmath__37[20]), .A0(N4905), .A1(N4925), .B0(N5085), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1136 (.Y(inst_cellmath__37[21]), .A0(N4905), .A1(N4972), .B0(N4916), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1137 (.Y(inst_cellmath__37[22]), .A0(N4905), .A1(N5017), .B0(N4965), .B1(N4953));
AOI22XL inst_cellmath__37_0_I3109 (.Y(inst_cellmath__37[23]), .A0(N4953), .A1(N5008), .B0(N4905), .B1(N5064));
AOI22XL inst_cellmath__37_0_I1139 (.Y(inst_cellmath__37[24]), .A0(N4905), .A1(N5114), .B0(N5057), .B1(N4953));
AOI22XL inst_cellmath__37_0_I3110 (.Y(inst_cellmath__37[25]), .A0(N4953), .A1(N5105), .B0(N4905), .B1(N4942));
AOI22XL inst_cellmath__37_0_I1141 (.Y(inst_cellmath__37[26]), .A0(N4905), .A1(N4993), .B0(N4935), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1142 (.Y(inst_cellmath__37[27]), .A0(N4905), .A1(N5036), .B0(N5029), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1143 (.Y(inst_cellmath__37[28]), .A0(N4905), .A1(N5085), .B0(N4907), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1144 (.Y(inst_cellmath__37[29]), .A0(N4905), .A1(N4916), .B0(N5003), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1145 (.Y(inst_cellmath__37[30]), .A0(N4905), .A1(N4965), .B0(N5097), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1146 (.Y(inst_cellmath__37[31]), .A0(N4905), .A1(N5008), .B0(N4977), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1147 (.Y(inst_cellmath__37[32]), .A0(N4905), .A1(N5057), .B0(N5070), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1148 (.Y(inst_cellmath__37[33]), .A0(N4905), .A1(N5105), .B0(N4948), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1149 (.Y(inst_cellmath__37[34]), .A0(N4905), .A1(N4935), .B0(N5041), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1150 (.Y(inst_cellmath__37[35]), .A0(N4905), .A1(N5029), .B0(N4922), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1151 (.Y(inst_cellmath__37[36]), .A0(N4905), .A1(N4907), .B0(N5014), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1152 (.Y(inst_cellmath__37[37]), .A0(N4905), .A1(N5003), .B0(N5111), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1153 (.Y(inst_cellmath__37[38]), .A0(N4905), .A1(N5097), .B0(N4990), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1154 (.Y(inst_cellmath__37[39]), .A0(N4905), .A1(N4977), .B0(N5081), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1155 (.Y(inst_cellmath__37[40]), .A0(N4905), .A1(N5070), .B0(N4960), .B1(N4953));
AOI22XL inst_cellmath__37_0_I1156 (.Y(inst_cellmath__37[41]), .A0(N4905), .A1(N4948), .B0(N5051), .B1(N4953));
NOR2XL inst_cellmath__37_0_I1164 (.Y(inst_cellmath__37[49]), .A(N4953), .B(N5051));
NOR2X1 inst_cellmath__33_49_24_I3205 (.Y(N5342), .A(inst_cellmath__31), .B(inst_cellmath__30));
AND2XL inst_cellmath__33_49_24_I1166 (.Y(inst_cellmath__33[24]), .A(N5342), .B(inst_cellmath__37[24]));
AND2XL inst_cellmath__33_49_24_I1167 (.Y(inst_cellmath__33[25]), .A(N5342), .B(inst_cellmath__37[25]));
AND2XL inst_cellmath__33_49_24_I1169 (.Y(inst_cellmath__33[27]), .A(N5342), .B(inst_cellmath__37[27]));
AND2XL inst_cellmath__33_49_24_I1171 (.Y(inst_cellmath__33[29]), .A(N5342), .B(inst_cellmath__37[29]));
AND2XL inst_cellmath__33_49_24_I1172 (.Y(inst_cellmath__33[30]), .A(N5342), .B(inst_cellmath__37[30]));
AND2XL inst_cellmath__33_49_24_I1173 (.Y(inst_cellmath__33[31]), .A(N5342), .B(inst_cellmath__37[31]));
AND2XL inst_cellmath__33_49_24_I1175 (.Y(inst_cellmath__33[33]), .A(N5342), .B(inst_cellmath__37[33]));
AND2XL inst_cellmath__33_49_24_I1177 (.Y(inst_cellmath__33[35]), .A(N5342), .B(inst_cellmath__37[35]));
AND2XL inst_cellmath__33_49_24_I1178 (.Y(inst_cellmath__33[36]), .A(N5342), .B(inst_cellmath__37[36]));
AND2XL inst_cellmath__33_49_24_I1179 (.Y(inst_cellmath__33[37]), .A(N5342), .B(inst_cellmath__37[37]));
AND2XL inst_cellmath__33_49_24_I1180 (.Y(inst_cellmath__33[38]), .A(N5342), .B(inst_cellmath__37[38]));
AND2XL inst_cellmath__33_49_24_I1181 (.Y(inst_cellmath__33[39]), .A(N5342), .B(inst_cellmath__37[39]));
AND2XL inst_cellmath__33_49_24_I1182 (.Y(inst_cellmath__33[40]), .A(N5342), .B(inst_cellmath__37[40]));
AND2XL inst_cellmath__33_49_24_I1183 (.Y(inst_cellmath__33[41]), .A(N5342), .B(inst_cellmath__37[41]));
NOR3BXL inst_cellmath__33_49_24_I3206 (.Y(inst_cellmath__33[42]), .AN(N5342), .B(N4953), .C(N5041));
NOR3BXL inst_cellmath__33_49_24_I3207 (.Y(inst_cellmath__33[43]), .AN(N5342), .B(N4953), .C(N4922));
NOR3BXL inst_cellmath__33_49_24_I3208 (.Y(inst_cellmath__33[44]), .AN(N5342), .B(N4953), .C(N5014));
NOR3BXL inst_cellmath__33_49_24_I3209 (.Y(inst_cellmath__33[45]), .AN(N5342), .B(N4953), .C(N5111));
NOR3BXL inst_cellmath__33_49_24_I3210 (.Y(inst_cellmath__33[46]), .AN(N5342), .B(N4953), .C(N4990));
NOR3BXL inst_cellmath__33_49_24_I3211 (.Y(inst_cellmath__33[47]), .AN(N5342), .B(N4953), .C(N5081));
NOR3BXL inst_cellmath__33_49_24_I3212 (.Y(inst_cellmath__33[48]), .AN(N5342), .B(N4953), .C(N4960));
NAND2XL inst_cellmath__33_49_24_I1191 (.Y(inst_cellmath__33[49]), .A(N5342), .B(inst_cellmath__37[49]));
NOR2XL inst_cellmath__42__22__I1192 (.Y(N5398), .A(inst_cellmath__30), .B(inst_cellmath__37[0]));
NOR2XL inst_cellmath__42__22__I1193 (.Y(N5408), .A(inst_cellmath__37[1]), .B(inst_cellmath__37[2]));
NAND2XL inst_cellmath__42__22__I1194 (.Y(N5419), .A(N5398), .B(N5408));
NOR2XL inst_cellmath__42__22__I1195 (.Y(N5428), .A(inst_cellmath__37[3]), .B(inst_cellmath__37[7]));
NOR2XL inst_cellmath__42__22__I1196 (.Y(N5437), .A(inst_cellmath__37[5]), .B(inst_cellmath__37[9]));
NOR2XL inst_cellmath__42__22__I1197 (.Y(N5402), .A(inst_cellmath__37[8]), .B(inst_cellmath__37[6]));
NOR2XL inst_cellmath__42__22__I1198 (.Y(N5411), .A(inst_cellmath__37[4]), .B(inst_cellmath__37[10]));
NOR2XL inst_cellmath__42__22__I1199 (.Y(N5431), .A(inst_cellmath__37[12]), .B(inst_cellmath__37[17]));
NOR2XL inst_cellmath__42__22__I1200 (.Y(N5416), .A(N5419), .B(inst_cellmath__37[19]));
NAND2XL inst_cellmath__42__22__I1201 (.Y(N5400), .A(N5428), .B(N5437));
NAND2XL inst_cellmath__42__22__I1202 (.Y(N5414), .A(N5402), .B(N5411));
NAND2XL inst_cellmath__42__22__I1203 (.Y(N5421), .A(N5416), .B(N5431));
NOR4X1 inst_cellmath__42__22__I1204 (.Y(N5407), .A(inst_cellmath__37[15]), .B(inst_cellmath__37[13]), .C(inst_cellmath__37[11]), .D(inst_cellmath__37[16]));
NOR3XL inst_cellmath__42__22__I1205 (.Y(N5404), .A(inst_cellmath__37[18]), .B(inst_cellmath__37[14]), .C(N5400));
NOR3XL inst_cellmath__42__22__I1206 (.Y(N5427), .A(inst_cellmath__37[23]), .B(inst_cellmath__37[22]), .C(N5414));
NOR3XL inst_cellmath__42__22__I1207 (.Y(N5397), .A(inst_cellmath__37[20]), .B(inst_cellmath__37[21]), .C(N5421));
NAND2XL inst_cellmath__42__22__I1208 (.Y(N5418), .A(N5407), .B(N5404));
NAND2XL inst_cellmath__42__22__I1209 (.Y(N5436), .A(N5427), .B(N5397));
OR2XL inst_cellmath__42__22__I1210 (.Y(N625), .A(N5418), .B(N5436));
NAND2BX1 cynw_cm_float_add2_ieee_I3067 (.Y(N8708), .AN(inst_cellmath__31), .B(N625));
INVX2 cynw_cm_float_add2_ieee_I3068 (.Y(inst_cellmath__42), .A(N8708));
INVX1 inst_cellmath__44_0_I1212 (.Y(N5465), .A(inst_cellmath__39[25]));
NOR3X4 inst_cellmath__44_0_I1213 (.Y(inst_cellmath__44), .A(N5465), .B(inst_cellmath__33[24]), .C(inst_cellmath__42));
MX2XL cynw_cm_float_add2_ieee_I1216 (.Y(N655), .A(a_man[0]), .B(b_man[0]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1217 (.Y(N656), .A(a_man[1]), .B(b_man[1]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1218 (.Y(N657), .A(a_man[2]), .B(b_man[2]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1219 (.Y(N658), .A(a_man[3]), .B(b_man[3]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1220 (.Y(N659), .A(a_man[4]), .B(b_man[4]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1221 (.Y(N660), .A(a_man[5]), .B(b_man[5]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1222 (.Y(N661), .A(a_man[6]), .B(b_man[6]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1223 (.Y(N662), .A(a_man[7]), .B(b_man[7]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1224 (.Y(N663), .A(a_man[8]), .B(b_man[8]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1225 (.Y(N664), .A(a_man[9]), .B(b_man[9]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1226 (.Y(N665), .A(a_man[10]), .B(b_man[10]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1227 (.Y(N666), .A(a_man[11]), .B(b_man[11]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1228 (.Y(N667), .A(a_man[12]), .B(b_man[12]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1229 (.Y(N668), .A(a_man[13]), .B(b_man[13]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1230 (.Y(N669), .A(a_man[14]), .B(b_man[14]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1231 (.Y(N670), .A(a_man[15]), .B(b_man[15]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1232 (.Y(N671), .A(a_man[16]), .B(b_man[16]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1233 (.Y(N672), .A(a_man[17]), .B(b_man[17]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1234 (.Y(N673), .A(a_man[18]), .B(b_man[18]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1235 (.Y(N674), .A(a_man[19]), .B(b_man[19]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1236 (.Y(N675), .A(a_man[20]), .B(b_man[20]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1237 (.Y(N676), .A(a_man[21]), .B(b_man[21]), .S0(N4832));
MX2XL cynw_cm_float_add2_ieee_I1238 (.Y(N677), .A(a_man[22]), .B(b_man[22]), .S0(N4832));
XNOR2X1 inst_cellmath__39__19__2mx_I1240 (.Y(inst_cellmath__39[0]), .A(inst_cellmath__33[25]), .B(N5465));
NAND2XL node_cs_const1_cs_ii_A_I3290 (.Y(N8861), .A(N5342), .B(inst_cellmath__37[26]));
XOR2XL node_cs_const1_cs_ii_A_I3291 (.Y(inst_cellmath__39[1]), .A(N5465), .B(N8861));
XNOR2X1 inst_cellmath__39__19__2mx_I1242 (.Y(inst_cellmath__39[2]), .A(inst_cellmath__33[27]), .B(N5465));
NAND2XL node_cs_const1_cs_ii_A_I3292 (.Y(N8868), .A(N5342), .B(inst_cellmath__37[28]));
XOR2XL node_cs_const1_cs_ii_A_I3293 (.Y(inst_cellmath__39[3]), .A(N5465), .B(N8868));
XNOR2X1 inst_cellmath__39__19__2mx_I1244 (.Y(inst_cellmath__39[4]), .A(inst_cellmath__33[29]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1245 (.Y(inst_cellmath__39[5]), .A(inst_cellmath__33[30]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1246 (.Y(inst_cellmath__39[6]), .A(inst_cellmath__33[31]), .B(N5465));
NAND2XL node_cs_const1_cs_ii_A_I3294 (.Y(N8875), .A(N5342), .B(inst_cellmath__37[32]));
XOR2XL node_cs_const1_cs_ii_A_I3295 (.Y(inst_cellmath__39[7]), .A(N5465), .B(N8875));
XNOR2X1 inst_cellmath__39__19__2mx_I1248 (.Y(inst_cellmath__39[8]), .A(inst_cellmath__33[33]), .B(N5465));
NAND2XL node_cs_const1_cs_ii_A_I3296 (.Y(N8882), .A(N5342), .B(inst_cellmath__37[34]));
XOR2XL node_cs_const1_cs_ii_A_I3297 (.Y(inst_cellmath__39[9]), .A(N5465), .B(N8882));
XNOR2X1 inst_cellmath__39__19__2mx_I1250 (.Y(inst_cellmath__39[10]), .A(inst_cellmath__33[35]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1251 (.Y(inst_cellmath__39[11]), .A(inst_cellmath__33[36]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1252 (.Y(inst_cellmath__39[12]), .A(inst_cellmath__33[37]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1253 (.Y(inst_cellmath__39[13]), .A(inst_cellmath__33[38]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1254 (.Y(inst_cellmath__39[14]), .A(inst_cellmath__33[39]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1255 (.Y(inst_cellmath__39[15]), .A(inst_cellmath__33[40]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1256 (.Y(inst_cellmath__39[16]), .A(inst_cellmath__33[41]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1257 (.Y(inst_cellmath__39[17]), .A(inst_cellmath__33[42]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1258 (.Y(inst_cellmath__39[18]), .A(inst_cellmath__33[43]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1259 (.Y(inst_cellmath__39[19]), .A(inst_cellmath__33[44]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1260 (.Y(inst_cellmath__39[20]), .A(inst_cellmath__33[45]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1261 (.Y(inst_cellmath__39[21]), .A(inst_cellmath__33[46]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1262 (.Y(inst_cellmath__39[22]), .A(inst_cellmath__33[47]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1263 (.Y(inst_cellmath__39[23]), .A(inst_cellmath__33[48]), .B(N5465));
XNOR2X1 inst_cellmath__39__19__2mx_I1264 (.Y(inst_cellmath__39[24]), .A(inst_cellmath__33[49]), .B(N5465));
NAND2X2 inst_cellmath__45_0_I1265 (.Y(N5725), .A(inst_cellmath__39[0]), .B(inst_cellmath__44));
NOR2XL inst_cellmath__45_0_I1266 (.Y(N5767), .A(N655), .B(inst_cellmath__39[1]));
XOR2XL inst_cellmath__45_0_I1267 (.Y(N5814), .A(N655), .B(inst_cellmath__39[1]));
NOR2XL inst_cellmath__45_0_I1268 (.Y(N5661), .A(N656), .B(inst_cellmath__39[2]));
XOR2XL inst_cellmath__45_0_I1269 (.Y(N5703), .A(N656), .B(inst_cellmath__39[2]));
NOR2XL inst_cellmath__45_0_I1270 (.Y(N5742), .A(N657), .B(inst_cellmath__39[3]));
XOR2XL inst_cellmath__45_0_I1271 (.Y(N5786), .A(N657), .B(inst_cellmath__39[3]));
NOR2XL inst_cellmath__45_0_I1272 (.Y(N5832), .A(N658), .B(inst_cellmath__39[4]));
XOR2XL inst_cellmath__45_0_I1273 (.Y(N5680), .A(N658), .B(inst_cellmath__39[4]));
NOR2XL inst_cellmath__45_0_I1274 (.Y(N5718), .A(N659), .B(inst_cellmath__39[5]));
XOR2XL inst_cellmath__45_0_I1275 (.Y(N5760), .A(N659), .B(inst_cellmath__39[5]));
NOR2XL inst_cellmath__45_0_I1276 (.Y(N5806), .A(N660), .B(inst_cellmath__39[6]));
XOR2XL inst_cellmath__45_0_I1277 (.Y(N5652), .A(N660), .B(inst_cellmath__39[6]));
NOR2XL inst_cellmath__45_0_I1278 (.Y(N5695), .A(N661), .B(inst_cellmath__39[7]));
XOR2XL inst_cellmath__45_0_I1279 (.Y(N5735), .A(N661), .B(inst_cellmath__39[7]));
NOR2XL inst_cellmath__45_0_I1280 (.Y(N5779), .A(N662), .B(inst_cellmath__39[8]));
XOR2XL inst_cellmath__45_0_I1281 (.Y(N5824), .A(N662), .B(inst_cellmath__39[8]));
NOR2XL inst_cellmath__45_0_I1282 (.Y(N5672), .A(N663), .B(inst_cellmath__39[9]));
XOR2XL inst_cellmath__45_0_I1283 (.Y(N5711), .A(N663), .B(inst_cellmath__39[9]));
NOR2XL inst_cellmath__45_0_I1284 (.Y(N5753), .A(N664), .B(inst_cellmath__39[10]));
XOR2XL inst_cellmath__45_0_I1285 (.Y(N5798), .A(N664), .B(inst_cellmath__39[10]));
NOR2XL inst_cellmath__45_0_I1286 (.Y(N5644), .A(N665), .B(inst_cellmath__39[11]));
XOR2XL inst_cellmath__45_0_I1287 (.Y(N5689), .A(N665), .B(inst_cellmath__39[11]));
NOR2XL inst_cellmath__45_0_I1288 (.Y(N5730), .A(N666), .B(inst_cellmath__39[12]));
XOR2XL inst_cellmath__45_0_I1289 (.Y(N5772), .A(N666), .B(inst_cellmath__39[12]));
NOR2XL inst_cellmath__45_0_I1290 (.Y(N5817), .A(N667), .B(inst_cellmath__39[13]));
XOR2XL inst_cellmath__45_0_I1291 (.Y(N5665), .A(N667), .B(inst_cellmath__39[13]));
NOR2XL inst_cellmath__45_0_I1292 (.Y(N5707), .A(N668), .B(inst_cellmath__39[14]));
XOR2XL inst_cellmath__45_0_I1293 (.Y(N5746), .A(N668), .B(inst_cellmath__39[14]));
NOR2XL inst_cellmath__45_0_I1294 (.Y(N5791), .A(N669), .B(inst_cellmath__39[15]));
XOR2XL inst_cellmath__45_0_I1295 (.Y(N5837), .A(N669), .B(inst_cellmath__39[15]));
NOR2XL inst_cellmath__45_0_I1296 (.Y(N5682), .A(N670), .B(inst_cellmath__39[16]));
XOR2XL inst_cellmath__45_0_I1297 (.Y(N5721), .A(N670), .B(inst_cellmath__39[16]));
NOR2XL inst_cellmath__45_0_I1298 (.Y(N5765), .A(N671), .B(inst_cellmath__39[17]));
XOR2XL inst_cellmath__45_0_I1299 (.Y(N5809), .A(N671), .B(inst_cellmath__39[17]));
NOR2XL inst_cellmath__45_0_I1300 (.Y(N5656), .A(N672), .B(inst_cellmath__39[18]));
XOR2XL inst_cellmath__45_0_I1301 (.Y(N5700), .A(N672), .B(inst_cellmath__39[18]));
NOR2XL inst_cellmath__45_0_I1302 (.Y(N5738), .A(N673), .B(inst_cellmath__39[19]));
XOR2XL inst_cellmath__45_0_I1303 (.Y(N5783), .A(N673), .B(inst_cellmath__39[19]));
NOR2XL inst_cellmath__45_0_I1304 (.Y(N5829), .A(N674), .B(inst_cellmath__39[20]));
XOR2XL inst_cellmath__45_0_I1305 (.Y(N5675), .A(N674), .B(inst_cellmath__39[20]));
NOR2XL inst_cellmath__45_0_I1306 (.Y(N5715), .A(N675), .B(inst_cellmath__39[21]));
XOR2XL inst_cellmath__45_0_I1307 (.Y(N5758), .A(N675), .B(inst_cellmath__39[21]));
NOR2XL inst_cellmath__45_0_I1308 (.Y(N5801), .A(N676), .B(inst_cellmath__39[22]));
XOR2XL inst_cellmath__45_0_I1309 (.Y(N5648), .A(N676), .B(inst_cellmath__39[22]));
NOR2XL inst_cellmath__45_0_I1310 (.Y(N5693), .A(N677), .B(inst_cellmath__39[23]));
XOR2XL inst_cellmath__45_0_I1311 (.Y(N5731), .A(N677), .B(inst_cellmath__39[23]));
AOI21X2 inst_cellmath__45_0_I1313 (.Y(N5668), .A0(N5814), .A1(N5725), .B0(N5767));
AOI21XL inst_cellmath__45_0_I1314 (.Y(N5749), .A0(N5786), .A1(N5661), .B0(N5742));
NAND2XL inst_cellmath__45_0_I1315 (.Y(N5792), .A(N5786), .B(N5703));
AOI21XL inst_cellmath__45_0_I1316 (.Y(N5839), .A0(N5760), .A1(N5832), .B0(N5718));
NAND2XL inst_cellmath__45_0_I1317 (.Y(N5686), .A(N5760), .B(N5680));
AOI21XL inst_cellmath__45_0_I1318 (.Y(N5723), .A0(N5735), .A1(N5806), .B0(N5695));
NAND2XL inst_cellmath__45_0_I1319 (.Y(N5766), .A(N5735), .B(N5652));
AOI21XL inst_cellmath__45_0_I1320 (.Y(N5813), .A0(N5711), .A1(N5779), .B0(N5672));
NAND2XL inst_cellmath__45_0_I1321 (.Y(N5660), .A(N5711), .B(N5824));
AOI21XL inst_cellmath__45_0_I1322 (.Y(N5702), .A0(N5689), .A1(N5753), .B0(N5644));
NAND2XL inst_cellmath__45_0_I1323 (.Y(N5741), .A(N5689), .B(N5798));
AOI21XL inst_cellmath__45_0_I1324 (.Y(N5785), .A0(N5665), .A1(N5730), .B0(N5817));
NAND2XL inst_cellmath__45_0_I1325 (.Y(N5831), .A(N5665), .B(N5772));
AOI21XL inst_cellmath__45_0_I1326 (.Y(N5679), .A0(N5837), .A1(N5707), .B0(N5791));
NAND2XL inst_cellmath__45_0_I1327 (.Y(N5717), .A(N5837), .B(N5746));
AOI21XL inst_cellmath__45_0_I1328 (.Y(N5759), .A0(N5809), .A1(N5682), .B0(N5765));
NAND2XL inst_cellmath__45_0_I1329 (.Y(N5805), .A(N5809), .B(N5721));
AOI21XL inst_cellmath__45_0_I1330 (.Y(N5651), .A0(N5783), .A1(N5656), .B0(N5738));
NAND2XL inst_cellmath__45_0_I1331 (.Y(N5694), .A(N5783), .B(N5700));
AOI21XL inst_cellmath__45_0_I1332 (.Y(N5734), .A0(N5758), .A1(N5829), .B0(N5715));
NAND2XL inst_cellmath__45_0_I1333 (.Y(N5778), .A(N5758), .B(N5675));
AOI21XL inst_cellmath__45_0_I1334 (.Y(N5823), .A0(N5731), .A1(N5801), .B0(N5693));
NAND2XL inst_cellmath__45_0_I1335 (.Y(N5671), .A(N5731), .B(N5648));
OAI21X2 inst_cellmath__45_0_I1336 (.Y(N5643), .A0(N5792), .A1(N5668), .B0(N5749));
OAI21XL inst_cellmath__45_0_I1337 (.Y(N5728), .A0(N5766), .A1(N5839), .B0(N5723));
NOR2XL inst_cellmath__45_0_I1338 (.Y(N5771), .A(N5766), .B(N5686));
OAI21XL inst_cellmath__45_0_I1339 (.Y(N5816), .A0(N5741), .A1(N5813), .B0(N5702));
NOR2XL inst_cellmath__45_0_I1340 (.Y(N5664), .A(N5741), .B(N5660));
OAI21XL inst_cellmath__45_0_I1341 (.Y(N5706), .A0(N5717), .A1(N5785), .B0(N5679));
NOR2XL inst_cellmath__45_0_I1342 (.Y(N5745), .A(N5717), .B(N5831));
OAI21XL inst_cellmath__45_0_I1343 (.Y(N5790), .A0(N5694), .A1(N5759), .B0(N5651));
NOR2XL inst_cellmath__45_0_I1344 (.Y(N5836), .A(N5694), .B(N5805));
AOI21X2 inst_cellmath__45_0_I1345 (.Y(N5763), .A0(N5771), .A1(N5643), .B0(N5728));
AOI21XL inst_cellmath__45_0_I1346 (.Y(N5655), .A0(N5745), .A1(N5816), .B0(N5706));
NAND2XL inst_cellmath__45_0_I1347 (.Y(N5698), .A(N5745), .B(N5664));
OAI21X2 inst_cellmath__45_0_I1348 (.Y(N5737), .A0(N5698), .A1(N5763), .B0(N5655));
INVXL inst_cellmath__45_0_I1349 (.Y(N5827), .A(N5664));
INVXL inst_cellmath__45_0_I1350 (.Y(N5674), .A(N5816));
OAI21XL inst_cellmath__45_0_I1351 (.Y(N5714), .A0(N5827), .A1(N5763), .B0(N5674));
INVXL inst_cellmath__45_0_I1352 (.Y(N5750), .A(N5737));
AOI21X2 inst_cellmath__45_0_I1353 (.Y(N5691), .A0(N5836), .A1(N5737), .B0(N5790));
INVXL inst_cellmath__45_0_I1354 (.Y(N5773), .A(N5686));
INVXL inst_cellmath__45_0_I1355 (.Y(N5820), .A(N5839));
AOI21XL inst_cellmath__45_0_I1356 (.Y(N5667), .A0(N5773), .A1(N5643), .B0(N5820));
INVXL inst_cellmath__45_0_I1357 (.Y(N5793), .A(N5763));
OAI21XL inst_cellmath__45_0_I1358 (.Y(N5838), .A0(N5660), .A1(N5763), .B0(N5813));
INVXL inst_cellmath__45_0_I1359 (.Y(N5840), .A(N5714));
INVXL inst_cellmath__45_0_I1360 (.Y(N5811), .A(N5831));
INVXL inst_cellmath__45_0_I1361 (.Y(N5659), .A(N5785));
AOI21XL inst_cellmath__45_0_I1362 (.Y(N5701), .A0(N5811), .A1(N5714), .B0(N5659));
INVXL inst_cellmath__45_0_I1363 (.Y(N5687), .A(N5750));
OAI21XL inst_cellmath__45_0_I1364 (.Y(N5677), .A0(N5805), .A1(N5750), .B0(N5759));
INVXL inst_cellmath__45_0_I1365 (.Y(N5724), .A(N5691));
OAI21X1 inst_cellmath__45_0_I1366 (.Y(N5650), .A0(N5778), .A1(N5691), .B0(N5734));
OA21X1 inst_cellmath__45_0_I1367 (.Y(N5777), .A0(N5671), .A1(N5734), .B0(N5823));
OAI31X1 inst_cellmath__45_0_I1368 (.Y(N5822), .A0(N5671), .A1(N5778), .A2(N5691), .B0(N5777));
INVXL inst_cellmath__45_0_I1369 (.Y(N5710), .A(N5703));
INVXL inst_cellmath__45_0_I1370 (.Y(N5752), .A(N5661));
OAI21XL inst_cellmath__45_0_I1371 (.Y(N5796), .A0(N5710), .A1(N5668), .B0(N5752));
AOI21XL inst_cellmath__45_0_I1372 (.Y(N5770), .A0(N5680), .A1(N5643), .B0(N5832));
INVXL inst_cellmath__45_0_I1373 (.Y(N5744), .A(N5652));
INVXL inst_cellmath__45_0_I1374 (.Y(N5788), .A(N5806));
OAI21XL inst_cellmath__45_0_I1375 (.Y(N5835), .A0(N5744), .A1(N5667), .B0(N5788));
AOI21XL inst_cellmath__45_0_I1376 (.Y(N5808), .A0(N5824), .A1(N5793), .B0(N5779));
AOI21XL inst_cellmath__45_0_I1377 (.Y(N5781), .A0(N5798), .A1(N5838), .B0(N5753));
INVXL inst_cellmath__45_0_I1378 (.Y(N5756), .A(N5772));
INVXL inst_cellmath__45_0_I1379 (.Y(N5800), .A(N5730));
OAI21XL inst_cellmath__45_0_I1380 (.Y(N5646), .A0(N5756), .A1(N5840), .B0(N5800));
INVXL inst_cellmath__45_0_I1381 (.Y(N5819), .A(N5746));
INVXL inst_cellmath__45_0_I1382 (.Y(N5666), .A(N5707));
OAI21XL inst_cellmath__45_0_I1383 (.Y(N5708), .A0(N5819), .A1(N5701), .B0(N5666));
AOI21XL inst_cellmath__45_0_I1384 (.Y(N5684), .A0(N5721), .A1(N5687), .B0(N5682));
AOI21XL inst_cellmath__45_0_I1385 (.Y(N5657), .A0(N5700), .A1(N5677), .B0(N5656));
AOI21XL inst_cellmath__45_0_I1386 (.Y(N5830), .A0(N5675), .A1(N5724), .B0(N5829));
AOI21XL inst_cellmath__45_0_I1387 (.Y(N5803), .A0(N5648), .A1(N5650), .B0(N5801));
NAND2XL inst_cellmath__45_0_I1388 (.Y(N5775), .A(inst_cellmath__39[24]), .B(N5822));
XOR2XL inst_cellmath__45_0_I1389 (.Y(inst_cellmath__45[0]), .A(inst_cellmath__39[0]), .B(inst_cellmath__44));
XNOR2X1 inst_cellmath__45_0_I1390 (.Y(inst_cellmath__45[1]), .A(N5725), .B(N5814));
XOR2XL inst_cellmath__45_0_I1391 (.Y(inst_cellmath__45[2]), .A(N5668), .B(N5703));
XNOR2X1 inst_cellmath__45_0_I1392 (.Y(inst_cellmath__45[3]), .A(N5796), .B(N5786));
XNOR2X1 inst_cellmath__45_0_I1393 (.Y(inst_cellmath__45[4]), .A(N5643), .B(N5680));
XOR2XL inst_cellmath__45_0_I1394 (.Y(inst_cellmath__45[5]), .A(N5770), .B(N5760));
XOR2XL inst_cellmath__45_0_I1395 (.Y(inst_cellmath__45[6]), .A(N5667), .B(N5652));
XNOR2X1 inst_cellmath__45_0_I1396 (.Y(inst_cellmath__45[7]), .A(N5835), .B(N5735));
XNOR2X1 inst_cellmath__45_0_I1397 (.Y(inst_cellmath__45[8]), .A(N5793), .B(N5824));
XOR2XL inst_cellmath__45_0_I1398 (.Y(inst_cellmath__45[9]), .A(N5808), .B(N5711));
XNOR2X1 inst_cellmath__45_0_I1399 (.Y(inst_cellmath__45[10]), .A(N5838), .B(N5798));
XOR2XL inst_cellmath__45_0_I1400 (.Y(inst_cellmath__45[11]), .A(N5781), .B(N5689));
XOR2XL inst_cellmath__45_0_I1401 (.Y(inst_cellmath__45[12]), .A(N5840), .B(N5772));
XNOR2X1 inst_cellmath__45_0_I1402 (.Y(inst_cellmath__45[13]), .A(N5646), .B(N5665));
XOR2XL inst_cellmath__45_0_I1403 (.Y(inst_cellmath__45[14]), .A(N5701), .B(N5746));
XNOR2X1 inst_cellmath__45_0_I1404 (.Y(inst_cellmath__45[15]), .A(N5708), .B(N5837));
XNOR2X1 inst_cellmath__45_0_I1405 (.Y(inst_cellmath__45[16]), .A(N5687), .B(N5721));
XOR2XL inst_cellmath__45_0_I1406 (.Y(inst_cellmath__45[17]), .A(N5684), .B(N5809));
XNOR2X1 inst_cellmath__45_0_I1407 (.Y(inst_cellmath__45[18]), .A(N5677), .B(N5700));
XOR2XL inst_cellmath__45_0_I1408 (.Y(inst_cellmath__45[19]), .A(N5657), .B(N5783));
XNOR2X1 inst_cellmath__45_0_I1409 (.Y(inst_cellmath__45[20]), .A(N5724), .B(N5675));
XOR2XL inst_cellmath__45_0_I1410 (.Y(inst_cellmath__45[21]), .A(N5830), .B(N5758));
XNOR2X1 inst_cellmath__45_0_I1411 (.Y(inst_cellmath__45[22]), .A(N5650), .B(N5648));
CLKXOR2X1 inst_cellmath__45_0_I1412 (.Y(inst_cellmath__45[23]), .A(N5803), .B(N5731));
XNOR2X1 inst_cellmath__45_0_I1413 (.Y(inst_cellmath__45[24]), .A(N5822), .B(inst_cellmath__39[24]));
XOR2XL inst_cellmath__45_0_I1414 (.Y(inst_cellmath__45[25]), .A(N5775), .B(inst_cellmath__39[25]));
NOR2BX1 inst_cellmath__49_0_I1415 (.Y(N6017), .AN(inst_cellmath__45[0]), .B(inst_cellmath__45[1]));
NOR2XL inst_cellmath__49_0_I1416 (.Y(N5996), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[0]));
NOR2BX1 inst_cellmath__49_0_I1417 (.Y(N6038), .AN(inst_cellmath__45[2]), .B(inst_cellmath__45[3]));
INVXL inst_cellmath__49_0_I1418 (.Y(N6057), .A(inst_cellmath__45[5]));
OAI21XL inst_cellmath__49_0_I1419 (.Y(N6079), .A0(inst_cellmath__45[4]), .A1(N6038), .B0(N6057));
NOR2XL inst_cellmath__49_0_I1420 (.Y(N6006), .A(inst_cellmath__45[3]), .B(inst_cellmath__45[2]));
NOR2XL inst_cellmath__49_0_I1421 (.Y(N6025), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[4]));
NOR2BX1 inst_cellmath__49_0_I1422 (.Y(N6067), .AN(inst_cellmath__45[6]), .B(inst_cellmath__45[7]));
INVXL inst_cellmath__49_0_I1423 (.Y(N6087), .A(inst_cellmath__45[9]));
OAI21XL inst_cellmath__49_0_I1424 (.Y(N6015), .A0(inst_cellmath__45[8]), .A1(N6067), .B0(N6087));
NOR2XL inst_cellmath__49_0_I1425 (.Y(N6033), .A(inst_cellmath__45[7]), .B(inst_cellmath__45[6]));
NOR2XL inst_cellmath__49_0_I1426 (.Y(N6052), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[8]));
NOR2BX1 inst_cellmath__49_0_I1427 (.Y(N6001), .AN(inst_cellmath__45[10]), .B(inst_cellmath__45[11]));
INVXL inst_cellmath__49_0_I1428 (.Y(N6021), .A(inst_cellmath__45[13]));
OAI21XL inst_cellmath__49_0_I1429 (.Y(N6043), .A0(inst_cellmath__45[12]), .A1(N6001), .B0(N6021));
NOR2XL inst_cellmath__49_0_I1430 (.Y(N6063), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[10]));
NOR2XL inst_cellmath__49_0_I1431 (.Y(N6083), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[12]));
NOR2BX1 inst_cellmath__49_0_I1432 (.Y(N6029), .AN(inst_cellmath__45[14]), .B(inst_cellmath__45[15]));
INVXL inst_cellmath__49_0_I1433 (.Y(N6050), .A(inst_cellmath__45[17]));
OAI21XL inst_cellmath__49_0_I1434 (.Y(N6071), .A0(inst_cellmath__45[16]), .A1(N6029), .B0(N6050));
NOR2X1 inst_cellmath__49_0_I1435 (.Y(N5998), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[14]));
NOR2X1 inst_cellmath__49_0_I1436 (.Y(N6019), .A(inst_cellmath__45[17]), .B(inst_cellmath__45[16]));
NOR2BX1 inst_cellmath__49_0_I1437 (.Y(N6058), .AN(inst_cellmath__45[18]), .B(inst_cellmath__45[19]));
INVXL inst_cellmath__49_0_I1438 (.Y(N6080), .A(inst_cellmath__45[21]));
OAI21XL inst_cellmath__49_0_I1439 (.Y(N6007), .A0(inst_cellmath__45[20]), .A1(N6058), .B0(N6080));
NOR2XL inst_cellmath__49_0_I1440 (.Y(N6026), .A(inst_cellmath__45[19]), .B(inst_cellmath__45[18]));
NOR2XL inst_cellmath__49_0_I1441 (.Y(N6047), .A(inst_cellmath__45[21]), .B(inst_cellmath__45[20]));
NOR2BX1 inst_cellmath__49_0_I1442 (.Y(N5993), .AN(inst_cellmath__45[22]), .B(inst_cellmath__45[23]));
INVXL inst_cellmath__49_0_I1443 (.Y(N6016), .A(inst_cellmath__45[25]));
OAI21XL inst_cellmath__49_0_I1444 (.Y(N6035), .A0(inst_cellmath__45[24]), .A1(N5993), .B0(N6016));
NOR2X1 inst_cellmath__49_0_I1445 (.Y(N6054), .A(inst_cellmath__45[23]), .B(inst_cellmath__45[22]));
NOR2X1 inst_cellmath__49_0_I1446 (.Y(N6076), .A(inst_cellmath__45[25]), .B(inst_cellmath__45[24]));
NAND2BXL inst_cellmath__49_0_I1447 (.Y(N6073), .AN(N6006), .B(N6025));
NAND2XL inst_cellmath__49_0_I1448 (.Y(N6041), .A(N6025), .B(N6006));
NAND2XL inst_cellmath__49_0_I1449 (.Y(N6060), .A(N6052), .B(N6033));
NAND2BXL inst_cellmath__49_0_I1450 (.Y(N6009), .AN(N6063), .B(N6083));
INVXL inst_cellmath__49_0_I1451 (.Y(N6028), .A(N6019));
AOI21XL inst_cellmath__49_0_I1452 (.Y(N6049), .A0(N5998), .A1(N6009), .B0(N6028));
NAND2XL inst_cellmath__49_0_I1453 (.Y(N6069), .A(N6083), .B(N6063));
NAND2X1 inst_cellmath__49_0_I1454 (.Y(N5995), .A(N6019), .B(N5998));
NAND2BXL inst_cellmath__49_0_I1455 (.Y(N6037), .AN(N6026), .B(N6047));
INVXL inst_cellmath__49_0_I1456 (.Y(N6056), .A(N6076));
AOI21XL inst_cellmath__49_0_I1457 (.Y(N6078), .A0(N6054), .A1(N6037), .B0(N6056));
NAND2XL inst_cellmath__49_0_I1458 (.Y(N6005), .A(N6047), .B(N6026));
NAND2X1 inst_cellmath__49_0_I1459 (.Y(N6024), .A(N6076), .B(N6054));
NAND2BXL inst_cellmath__49_0_I1460 (.Y(N6014), .AN(N6060), .B(N6041));
NOR2XL inst_cellmath__49_0_I1461 (.Y(N6000), .A(N6060), .B(N6041));
NOR2BX1 inst_cellmath__49_0_I1462 (.Y(N6042), .AN(N6069), .B(N5995));
INVXL inst_cellmath__49_0_I1463 (.Y(N6062), .A(N6024));
OAI21XL inst_cellmath__49_0_I1464 (.Y(N6082), .A0(N6005), .A1(N6042), .B0(N6062));
NOR2X1 inst_cellmath__49_0_I1465 (.Y(N6011), .A(N5995), .B(N6069));
NOR2X1 inst_cellmath__49_0_I1466 (.Y(N6061), .A(N6024), .B(N6005));
NAND2BXL inst_cellmath__49_0_I1467 (.Y(N6070), .AN(N5996), .B(N6000));
INVXL inst_cellmath__49_0_I1468 (.Y(N5997), .A(N6061));
NAND2XL inst_cellmath__49_0_I1470 (.Y(N6039), .A(N6000), .B(N5996));
NAND2X1 inst_cellmath__49_0_I1471 (.Y(N6010), .A(N6011), .B(N6061));
NOR2XL inst_cellmath__49_0_I1473 (.Y(inst_cellmath__49[5]), .A(N6010), .B(N6039));
OAI2BB1X1 inst_cellmath__49_0_I1475 (.Y(N6065), .A0N(N6033), .A1N(N6073), .B0(N6052));
AOI21XL inst_cellmath__49_0_I1476 (.Y(N6031), .A0(N6061), .A1(N6049), .B0(N6078));
OAI21X2 inst_cellmath__49_0_I1477 (.Y(inst_cellmath__49[1]), .A0(N6010), .A1(N6065), .B0(N6031));
OAI21XL inst_cellmath__49_0_I1478 (.Y(N6004), .A0(N6060), .A1(N6079), .B0(N6015));
OAI21XL inst_cellmath__49_0_I1479 (.Y(N6046), .A0(N5995), .A1(N6043), .B0(N6071));
OAI21XL inst_cellmath__49_0_I1480 (.Y(N6086), .A0(N6024), .A1(N6007), .B0(N6035));
AOI21XL inst_cellmath__49_0_I1481 (.Y(N6032), .A0(N6000), .A1(N6017), .B0(N6004));
AOI21XL inst_cellmath__49_0_I1482 (.Y(N6074), .A0(N6061), .A1(N6046), .B0(N6086));
OAI21X2 inst_cellmath__49_0_I1483 (.Y(inst_cellmath__49[0]), .A0(N6010), .A1(N6032), .B0(N6074));
OR2XL cmp_A_I7972 (.Y(N13895), .A(a_sign), .B(b_sign));
AO22XL cmp_A_I7973 (.Y(N645), .A0(N13895), .A1(inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL cynw_cm_float_add2_ieee_I1489 (.Y(inst_cellmath__66), .A(inst_cellmath__11), .B(N645), .C(inst_cellmath__16));
NOR2BX1 inst_cellmath__64__48__2WWMM_I1490 (.Y(N6212), .AN(inst_cellmath__18), .B(inst_cellmath__13));
AOI22XL inst_cellmath__64__48__2WWMM_I1491 (.Y(N6233), .A0(a_sign), .A1(inst_cellmath__13), .B0(N6212), .B1(b_sign));
AO22XL inst_cellmath__64__48__2WWMM_I1492 (.Y(inst_cellmath__64[0]), .A0(inst_cellmath__13), .A1(a_man[0]), .B0(N6212), .B1(b_man[0]));
AO22XL inst_cellmath__64__48__2WWMM_I1493 (.Y(inst_cellmath__64[1]), .A0(inst_cellmath__13), .A1(a_man[1]), .B0(N6212), .B1(b_man[1]));
AO22XL inst_cellmath__64__48__2WWMM_I1494 (.Y(inst_cellmath__64[2]), .A0(inst_cellmath__13), .A1(a_man[2]), .B0(N6212), .B1(b_man[2]));
AO22XL inst_cellmath__64__48__2WWMM_I1495 (.Y(inst_cellmath__64[3]), .A0(inst_cellmath__13), .A1(a_man[3]), .B0(N6212), .B1(b_man[3]));
AO22XL inst_cellmath__64__48__2WWMM_I1496 (.Y(inst_cellmath__64[4]), .A0(inst_cellmath__13), .A1(a_man[4]), .B0(N6212), .B1(b_man[4]));
AO22XL inst_cellmath__64__48__2WWMM_I1497 (.Y(inst_cellmath__64[5]), .A0(inst_cellmath__13), .A1(a_man[5]), .B0(N6212), .B1(b_man[5]));
AO22XL inst_cellmath__64__48__2WWMM_I1498 (.Y(inst_cellmath__64[6]), .A0(inst_cellmath__13), .A1(a_man[6]), .B0(N6212), .B1(b_man[6]));
AO22XL inst_cellmath__64__48__2WWMM_I1499 (.Y(inst_cellmath__64[7]), .A0(inst_cellmath__13), .A1(a_man[7]), .B0(N6212), .B1(b_man[7]));
AO22XL inst_cellmath__64__48__2WWMM_I1500 (.Y(inst_cellmath__64[8]), .A0(inst_cellmath__13), .A1(a_man[8]), .B0(N6212), .B1(b_man[8]));
AO22XL inst_cellmath__64__48__2WWMM_I1501 (.Y(inst_cellmath__64[9]), .A0(inst_cellmath__13), .A1(a_man[9]), .B0(N6212), .B1(b_man[9]));
AO22XL inst_cellmath__64__48__2WWMM_I1502 (.Y(inst_cellmath__64[10]), .A0(inst_cellmath__13), .A1(a_man[10]), .B0(N6212), .B1(b_man[10]));
AO22XL inst_cellmath__64__48__2WWMM_I1503 (.Y(inst_cellmath__64[11]), .A0(inst_cellmath__13), .A1(a_man[11]), .B0(N6212), .B1(b_man[11]));
AO22XL inst_cellmath__64__48__2WWMM_I1504 (.Y(inst_cellmath__64[12]), .A0(inst_cellmath__13), .A1(a_man[12]), .B0(N6212), .B1(b_man[12]));
AO22XL inst_cellmath__64__48__2WWMM_I1505 (.Y(inst_cellmath__64[13]), .A0(inst_cellmath__13), .A1(a_man[13]), .B0(N6212), .B1(b_man[13]));
AO22XL inst_cellmath__64__48__2WWMM_I1506 (.Y(inst_cellmath__64[14]), .A0(inst_cellmath__13), .A1(a_man[14]), .B0(N6212), .B1(b_man[14]));
AO22XL inst_cellmath__64__48__2WWMM_I1507 (.Y(inst_cellmath__64[15]), .A0(inst_cellmath__13), .A1(a_man[15]), .B0(N6212), .B1(b_man[15]));
AO22XL inst_cellmath__64__48__2WWMM_I1508 (.Y(inst_cellmath__64[16]), .A0(inst_cellmath__13), .A1(a_man[16]), .B0(N6212), .B1(b_man[16]));
AO22XL inst_cellmath__64__48__2WWMM_I1509 (.Y(inst_cellmath__64[17]), .A0(inst_cellmath__13), .A1(a_man[17]), .B0(N6212), .B1(b_man[17]));
AO22XL inst_cellmath__64__48__2WWMM_I1510 (.Y(inst_cellmath__64[18]), .A0(inst_cellmath__13), .A1(a_man[18]), .B0(N6212), .B1(b_man[18]));
AO22XL inst_cellmath__64__48__2WWMM_I1511 (.Y(inst_cellmath__64[19]), .A0(inst_cellmath__13), .A1(a_man[19]), .B0(N6212), .B1(b_man[19]));
AO22XL inst_cellmath__64__48__2WWMM_I1512 (.Y(inst_cellmath__64[20]), .A0(inst_cellmath__13), .A1(a_man[20]), .B0(N6212), .B1(b_man[20]));
AO22XL inst_cellmath__64__48__2WWMM_I1513 (.Y(inst_cellmath__64[21]), .A0(inst_cellmath__13), .A1(a_man[21]), .B0(N6212), .B1(b_man[21]));
OAI21XL inst_cellmath__64__48__2WWMM_I1514 (.Y(N710), .A0(inst_cellmath__18), .A1(inst_cellmath__13), .B0(N6233));
MX2XL inst_cellmath__67_0_I1515 (.Y(N6282), .A(inst_cellmath__66), .B(N710), .S0(inst_cellmath__63));
NOR2XL inst_cellmath__67_0_I1516 (.Y(N6291), .A(inst_cellmath__63), .B(N706));
MX2XL inst_cellmath__67_0_I7942 (.Y(N6285), .A(inst_cellmath__48), .B(inst_cellmath__6), .S0(inst_cellmath__49[5]));
MX2XL inst_cellmath__67_0_I1518 (.Y(x[31]), .A(N6282), .B(N6285), .S0(N6291));
AO21X1 inst_cellmath__50_0_I3221 (.Y(N6439), .A0(N6011), .A1(N6070), .B0(N5997));
INVX1 inst_cellmath__50_0_I3169 (.Y(N8804), .A(N6439));
INVX1 inst_cellmath__50_0_I3174 (.Y(N8809), .A(N8804));
INVX1 inst_cellmath__50_0_I3173 (.Y(N8808), .A(N8804));
INVXL inst_cellmath__50_0_I3171 (.Y(N8806), .A(N8804));
AND2X1 inst_cellmath__50_0_I1520 (.Y(N6312), .A(inst_cellmath__45[0]), .B(N6439));
AND2XL inst_cellmath__50_0_I1521 (.Y(N6383), .A(inst_cellmath__45[1]), .B(N8809));
CLKAND2X2 inst_cellmath__50_0_I1522 (.Y(N6454), .A(N8809), .B(inst_cellmath__45[2]));
AND2XL inst_cellmath__50_0_I1523 (.Y(N6361), .A(N8809), .B(inst_cellmath__45[3]));
AND2XL inst_cellmath__50_0_I1524 (.Y(N6432), .A(N8809), .B(inst_cellmath__45[4]));
AND2XL inst_cellmath__50_0_I1525 (.Y(N6341), .A(N8808), .B(inst_cellmath__45[5]));
AND2XL inst_cellmath__50_0_I1526 (.Y(N6411), .A(N8808), .B(inst_cellmath__45[6]));
AND2XL inst_cellmath__50_0_I1527 (.Y(N6321), .A(N8808), .B(inst_cellmath__45[7]));
MX2XL inst_cellmath__50_0_I1528 (.Y(N6392), .A(inst_cellmath__45[0]), .B(inst_cellmath__45[8]), .S0(N8808));
MX2XL inst_cellmath__50_0_I1529 (.Y(N6427), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[9]), .S0(N8808));
MX2XL inst_cellmath__50_0_I1530 (.Y(N6297), .A(inst_cellmath__45[2]), .B(inst_cellmath__45[10]), .S0(N8808));
MX2XL inst_cellmath__50_0_I1531 (.Y(N6334), .A(inst_cellmath__45[3]), .B(inst_cellmath__45[11]), .S0(N8808));
MX2XL inst_cellmath__50_0_I1532 (.Y(N6371), .A(inst_cellmath__45[4]), .B(inst_cellmath__45[12]), .S0(N8808));
MX2XL inst_cellmath__50_0_I1533 (.Y(N6405), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[13]), .S0(N8808));
MX2XL inst_cellmath__50_0_I1534 (.Y(N6441), .A(inst_cellmath__45[6]), .B(inst_cellmath__45[14]), .S0(N8808));
MX2XL inst_cellmath__50_0_I1535 (.Y(N6315), .A(inst_cellmath__45[7]), .B(inst_cellmath__45[15]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1536 (.Y(N6349), .A(inst_cellmath__45[8]), .B(inst_cellmath__45[16]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1537 (.Y(N6386), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[17]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1538 (.Y(N6420), .A(inst_cellmath__45[10]), .B(inst_cellmath__45[18]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1539 (.Y(N6457), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[19]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1540 (.Y(N6328), .A(inst_cellmath__45[12]), .B(inst_cellmath__45[20]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1541 (.Y(N6365), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[21]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1542 (.Y(N6400), .A(inst_cellmath__45[14]), .B(inst_cellmath__45[22]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1543 (.Y(N6436), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[23]), .S0(N8806));
MX2XL inst_cellmath__50_0_I1544 (.Y(N6307), .A(inst_cellmath__45[16]), .B(inst_cellmath__45[24]), .S0(N8806));
NAND2BX2 inst_cellmath__50_0_I3222 (.Y(N6311), .AN(N6010), .B(N6039));
INVXL inst_cellmath__50_0_I1546 (.Y(N6347), .A(N6311));
NAND2X1 inst_cellmath__50_0_I1547 (.Y(N6303), .A(N6311), .B(N6312));
NAND2X1 inst_cellmath__50_0_I1548 (.Y(N6377), .A(N6311), .B(N6383));
NAND2X1 inst_cellmath__50_0_I1549 (.Y(N6447), .A(N6311), .B(N6454));
NAND2XL inst_cellmath__50_0_I1550 (.Y(N6355), .A(N6361), .B(N6311));
NAND2XL inst_cellmath__50_0_I1551 (.Y(N6426), .A(N6432), .B(N6311));
NAND2XL inst_cellmath__50_0_I1552 (.Y(N6333), .A(N6341), .B(N6311));
NAND2XL inst_cellmath__50_0_I1553 (.Y(N6404), .A(N6411), .B(N6311));
NAND2XL inst_cellmath__50_0_I1554 (.Y(N6314), .A(N6321), .B(N6311));
NAND2XL inst_cellmath__50_0_I1555 (.Y(N6385), .A(N6392), .B(N6311));
NAND2XL inst_cellmath__50_0_I1556 (.Y(N6456), .A(N6427), .B(N6311));
NAND2XL inst_cellmath__50_0_I1557 (.Y(N6364), .A(N6297), .B(N6311));
NAND2XL inst_cellmath__50_0_I1558 (.Y(N6435), .A(N6334), .B(N6311));
NAND2XL inst_cellmath__50_0_I1559 (.Y(N6344), .A(N6371), .B(N6311));
NAND2XL inst_cellmath__50_0_I1560 (.Y(N6414), .A(N6405), .B(N6311));
NAND2XL inst_cellmath__50_0_I1561 (.Y(N6324), .A(N6441), .B(N6311));
NAND2XL inst_cellmath__50_0_I1562 (.Y(N6395), .A(N6315), .B(N6311));
AOI22XL inst_cellmath__50_0_I1563 (.Y(N6300), .A0(N6347), .A1(N6312), .B0(N6349), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1564 (.Y(N6337), .A0(N6347), .A1(N6383), .B0(N6386), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1565 (.Y(N6374), .A0(N6347), .A1(N6454), .B0(N6420), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1566 (.Y(N6408), .A0(N6347), .A1(N6361), .B0(N6457), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1567 (.Y(N6444), .A0(N6347), .A1(N6432), .B0(N6328), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1568 (.Y(N6318), .A0(N6347), .A1(N6341), .B0(N6365), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1569 (.Y(N6352), .A0(N6347), .A1(N6411), .B0(N6400), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1570 (.Y(N6389), .A0(N6347), .A1(N6321), .B0(N6436), .B1(N6311));
AOI22XL inst_cellmath__50_0_I1571 (.Y(N6423), .A0(N6347), .A1(N6392), .B0(N6307), .B1(N6311));
INVX2 inst_cellmath__50_0_I1572 (.Y(N6416), .A(inst_cellmath__49[0]));
INVX1 inst_cellmath__50_0_I1573 (.Y(N6452), .A(N6416));
INVX1 inst_cellmath__50_0_I3177 (.Y(N8812), .A(N6452));
INVX1 inst_cellmath__50_0_I3182 (.Y(N8817), .A(N8812));
INVXL inst_cellmath__50_0_I3181 (.Y(N8816), .A(N8812));
INVXL inst_cellmath__50_0_I3179 (.Y(N8814), .A(N8812));
NOR2XL inst_cellmath__50_0_I1574 (.Y(N6419), .A(N6452), .B(N6303));
AOI22XL inst_cellmath__50_0_I1575 (.Y(N6362), .A0(N6416), .A1(N6377), .B0(N6303), .B1(N8814));
AOI22X2 inst_cellmath__50_0_I1576 (.Y(N6398), .A0(N6416), .A1(N6447), .B0(N6377), .B1(N8817));
AOI22XL inst_cellmath__50_0_I1577 (.Y(N6434), .A0(N6416), .A1(N6355), .B0(N6447), .B1(N8817));
AOI22XL inst_cellmath__50_0_I1578 (.Y(N6306), .A0(N6416), .A1(N6426), .B0(N6355), .B1(N8817));
AOI22XL inst_cellmath__50_0_I1579 (.Y(N6343), .A0(N6416), .A1(N6333), .B0(N6426), .B1(N8817));
AOI22XL inst_cellmath__50_0_I1580 (.Y(N6379), .A0(N6416), .A1(N6404), .B0(N6333), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1581 (.Y(N6412), .A0(N6416), .A1(N6314), .B0(N6404), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1582 (.Y(N6448), .A0(N6416), .A1(N6385), .B0(N6314), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1583 (.Y(N6323), .A0(N6416), .A1(N6456), .B0(N6385), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1584 (.Y(N6357), .A0(N6416), .A1(N6364), .B0(N6456), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1585 (.Y(N6394), .A0(N6416), .A1(N6435), .B0(N6364), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1586 (.Y(N6429), .A0(N6416), .A1(N6344), .B0(N6435), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1587 (.Y(N6298), .A0(N6416), .A1(N6414), .B0(N6344), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1588 (.Y(N6335), .A0(N6416), .A1(N6324), .B0(N6414), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1589 (.Y(N6373), .A0(N6416), .A1(N6395), .B0(N6324), .B1(N8816));
AOI22XL inst_cellmath__50_0_I1590 (.Y(N6407), .A0(N6416), .A1(N6300), .B0(N6395), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1591 (.Y(N6443), .A0(N6416), .A1(N6337), .B0(N6300), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1592 (.Y(N6317), .A0(N6416), .A1(N6374), .B0(N6337), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1593 (.Y(N6350), .A0(N6416), .A1(N6408), .B0(N6374), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1594 (.Y(N6387), .A0(N6416), .A1(N6444), .B0(N6408), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1595 (.Y(N6422), .A0(N6416), .A1(N6318), .B0(N6444), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1596 (.Y(N6459), .A0(N6416), .A1(N6352), .B0(N6318), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1597 (.Y(N6330), .A0(N6416), .A1(N6389), .B0(N6352), .B1(N8814));
AOI22XL inst_cellmath__50_0_I1598 (.Y(N6367), .A0(N6416), .A1(N6423), .B0(N6389), .B1(N8814));
OA21X1 inst_cellmath__50_0_I3223 (.Y(N6360), .A0(N6014), .A1(N6010), .B0(N6082));
INVX1 inst_cellmath__50_0_I1600 (.Y(N6397), .A(N6360));
NAND2X1 inst_cellmath__50_0_I1601 (.Y(N6308), .A(N6419), .B(N6360));
NAND2XL inst_cellmath__50_0_I1602 (.Y(N6380), .A(N6362), .B(N6360));
NAND2X1 inst_cellmath__50_0_I1603 (.Y(N6450), .A(N6360), .B(N6398));
NAND2XL inst_cellmath__50_0_I1604 (.Y(N6358), .A(N6434), .B(N6360));
AOI22XL inst_cellmath__50_0_I1605 (.Y(N6430), .A0(N6397), .A1(N6419), .B0(N6306), .B1(N6360));
AOI22XL inst_cellmath__50_0_I3118 (.Y(N6301), .A0(N6343), .A1(N6360), .B0(N6397), .B1(N6362));
AOI22XL inst_cellmath__50_0_I1607 (.Y(N6338), .A0(N6397), .A1(N6398), .B0(N6379), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1608 (.Y(N6375), .A0(N6397), .A1(N6434), .B0(N6412), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1609 (.Y(N6409), .A0(N6397), .A1(N6306), .B0(N6448), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1610 (.Y(N6445), .A0(N6397), .A1(N6343), .B0(N6323), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1611 (.Y(N6319), .A0(N6397), .A1(N6379), .B0(N6357), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1612 (.Y(N6353), .A0(N6397), .A1(N6412), .B0(N6394), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1613 (.Y(N6390), .A0(N6397), .A1(N6448), .B0(N6429), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1614 (.Y(N6424), .A0(N6397), .A1(N6323), .B0(N6298), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1615 (.Y(N6460), .A0(N6397), .A1(N6357), .B0(N6335), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1616 (.Y(N6331), .A0(N6397), .A1(N6394), .B0(N6373), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1617 (.Y(N6368), .A0(N6397), .A1(N6429), .B0(N6407), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1618 (.Y(N6402), .A0(N6397), .A1(N6298), .B0(N6443), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1619 (.Y(N6438), .A0(N6397), .A1(N6335), .B0(N6317), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1620 (.Y(N6310), .A0(N6397), .A1(N6373), .B0(N6350), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1621 (.Y(N6346), .A0(N6397), .A1(N6407), .B0(N6387), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1622 (.Y(N6382), .A0(N6397), .A1(N6443), .B0(N6422), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1623 (.Y(N6417), .A0(N6397), .A1(N6317), .B0(N6459), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1624 (.Y(N6453), .A0(N6397), .A1(N6350), .B0(N6330), .B1(N6360));
AOI22XL inst_cellmath__50_0_I1625 (.Y(N6326), .A0(N6397), .A1(N6387), .B0(N6367), .B1(N6360));
INVXL inst_cellmath__50_0_I3189 (.Y(N8824), .A(inst_cellmath__49[1]));
INVXL inst_cellmath__50_0_I3185 (.Y(N8820), .A(inst_cellmath__49[1]));
NOR2XL inst_cellmath__50_0_I1629 (.Y(inst_cellmath__50[1]), .A(inst_cellmath__49[1]), .B(N6380));
AOI22XL inst_cellmath__50_0_I3087 (.Y(N8772), .A0(N8820), .A1(N6450), .B0(N6308), .B1(inst_cellmath__49[1]));
INVXL inst_cellmath__50_0_I3088 (.Y(inst_cellmath__50[2]), .A(N8772));
AOI22XL inst_cellmath__50_0_I1631 (.Y(inst_cellmath__50[3]), .A0(N8824), .A1(N6358), .B0(N6380), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1632 (.Y(inst_cellmath__50[4]), .A0(N8824), .A1(N6430), .B0(N6450), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I3119 (.Y(inst_cellmath__50[5]), .A0(inst_cellmath__49[1]), .A1(N6358), .B0(N8820), .B1(N6301));
AOI22XL inst_cellmath__50_0_I1634 (.Y(inst_cellmath__50[6]), .A0(N8824), .A1(N6338), .B0(N6430), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I3120 (.Y(inst_cellmath__50[7]), .A0(inst_cellmath__49[1]), .A1(N6301), .B0(N8820), .B1(N6375));
AOI22XL inst_cellmath__50_0_I1636 (.Y(inst_cellmath__50[8]), .A0(N8824), .A1(N6409), .B0(N6338), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1637 (.Y(inst_cellmath__50[9]), .A0(N8824), .A1(N6445), .B0(N6375), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1638 (.Y(inst_cellmath__50[10]), .A0(N8824), .A1(N6319), .B0(N6409), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1639 (.Y(inst_cellmath__50[11]), .A0(N8824), .A1(N6353), .B0(N6445), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1640 (.Y(inst_cellmath__50[12]), .A0(N8824), .A1(N6390), .B0(N6319), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1641 (.Y(inst_cellmath__50[13]), .A0(N8824), .A1(N6424), .B0(N6353), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1642 (.Y(inst_cellmath__50[14]), .A0(N8824), .A1(N6460), .B0(N6390), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1643 (.Y(inst_cellmath__50[15]), .A0(N8824), .A1(N6331), .B0(N6424), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1644 (.Y(inst_cellmath__50[16]), .A0(N8824), .A1(N6368), .B0(N6460), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1645 (.Y(inst_cellmath__50[17]), .A0(N8824), .A1(N6402), .B0(N6331), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1646 (.Y(inst_cellmath__50[18]), .A0(N8824), .A1(N6438), .B0(N6368), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1647 (.Y(inst_cellmath__50[19]), .A0(N8824), .A1(N6310), .B0(N6402), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1648 (.Y(inst_cellmath__50[20]), .A0(N8820), .A1(N6346), .B0(N6438), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1649 (.Y(inst_cellmath__50[21]), .A0(N8820), .A1(N6382), .B0(N6310), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1650 (.Y(inst_cellmath__50[22]), .A0(N8820), .A1(N6417), .B0(N6346), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1651 (.Y(inst_cellmath__50[23]), .A0(N8820), .A1(N6453), .B0(N6382), .B1(inst_cellmath__49[1]));
AOI22XL inst_cellmath__50_0_I1652 (.Y(inst_cellmath__50[24]), .A0(N8820), .A1(N6326), .B0(N6417), .B1(inst_cellmath__49[1]));
XNOR2X1 cynw_cm_float_add2_ieee_I1653 (.Y(N626), .A(inst_cellmath__33[24]), .B(inst_cellmath__42));
OR2XL cynw_cm_float_add2_ieee_I1655 (.Y(N627), .A(inst_cellmath__30), .B(N626));
OR2XL cynw_cm_float_add2_ieee_I1656 (.Y(N628), .A(inst_cellmath__33[24]), .B(inst_cellmath__42));
OAI2BB1X1 cynw_cm_float_add2_ieee_I3225 (.Y(N630), .A0N(inst_cellmath__30), .A1N(N628), .B0(N627));
MX2XL cynw_cm_float_add2_ieee_I1659 (.Y(inst_cellmath__43), .A(inst_cellmath__33[24]), .B(N630), .S0(inst_cellmath__39[25]));
MXI2XL cynw_cm_float_add2_ieee_I1660 (.Y(inst_cellmath__53), .A(inst_cellmath__50[1]), .B(inst_cellmath__43), .S0(inst_cellmath__49[1]));
NOR3BXL cynw_cm_float_add2_ieee_I1661 (.Y(inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
NOR2BX1 cynw_cm_float_add2_ieee_I3226 (.Y(N635), .AN(inst_cellmath__5), .B(inst_cellmath__48));
AND2XL cynw_cm_float_add2_ieee_I1664 (.Y(N634), .A(inst_cellmath__6), .B(inst_cellmath__48));
NOR3BXL cynw_cm_float_add2_ieee_I1665 (.Y(inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3XL cynw_cm_float_add2_ieee_I1666 (.Y(inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
NOR2XL inst_cellmath__54__33__I1667 (.Y(N6655), .A(inst_cellmath__42), .B(inst_cellmath__43));
OAI21XL inst_cellmath__54__33__I3228 (.Y(N631), .A0(inst_cellmath__49[1]), .A1(N6308), .B0(N6655));
MXI2XL cynw_cm_float_add2_ieee_I3149 (.Y(inst_cellmath__54), .A(N631), .B(inst_cellmath__42), .S0(inst_cellmath__49[1]));
NAND2XL cynw_cm_float_add2_ieee_I1670 (.Y(N632), .A(inst_cellmath__50[2]), .B(inst_cellmath__54));
AND2XL cynw_cm_float_add2_ieee_I1671 (.Y(N633), .A(inst_cellmath__4), .B(N632));
NOR4X1 cynw_cm_float_add2_ieee_I1672 (.Y(N636), .A(inst_cellmath__8), .B(N635), .C(N634), .D(N633));
NOR2XL cynw_cm_float_add2_ieee_I1674 (.Y(N638), .A(N635), .B(N634));
NOR2XL cynw_cm_float_add2_ieee_I1675 (.Y(N639), .A(N638), .B(inst_cellmath__54));
AOI2BB1XL cynw_cm_float_add2_ieee_I3122 (.Y(inst_cellmath__55), .A0N(inst_cellmath__53), .A1N(N636), .B0(N639));
OR2X1 inst_cellmath__57_0_I1677 (.Y(N6776), .A(inst_cellmath__55), .B(inst_cellmath__50[2]));
NAND2XL inst_cellmath__57_0_I1678 (.Y(N6719), .A(inst_cellmath__50[6]), .B(inst_cellmath__50[5]));
NAND2XL inst_cellmath__57_0_I1679 (.Y(N6709), .A(inst_cellmath__50[10]), .B(inst_cellmath__50[9]));
NAND2XL inst_cellmath__57_0_I1680 (.Y(N6727), .A(inst_cellmath__50[14]), .B(inst_cellmath__50[13]));
NAND2XL inst_cellmath__57_0_I1681 (.Y(N6767), .A(inst_cellmath__50[18]), .B(inst_cellmath__50[17]));
NAND2XL inst_cellmath__57_0_I1682 (.Y(N6769), .A(inst_cellmath__50[4]), .B(inst_cellmath__50[3]));
NOR2X2 inst_cellmath__57_0_I1683 (.Y(N6731), .A(N6776), .B(N6769));
NAND2XL inst_cellmath__57_0_I1684 (.Y(N6734), .A(inst_cellmath__50[12]), .B(inst_cellmath__50[11]));
NOR2X1 inst_cellmath__57_0_I1685 (.Y(N6751), .A(N6709), .B(N6734));
NAND4BX2 inst_cellmath__57_0_I1686 (.Y(N6759), .AN(N6719), .B(inst_cellmath__50[7]), .C(inst_cellmath__50[8]), .D(N6731));
NAND4BX1 inst_cellmath__57_0_I1687 (.Y(N6749), .AN(N6727), .B(inst_cellmath__50[15]), .C(inst_cellmath__50[16]), .D(N6751));
NOR2X1 inst_cellmath__57_0_I1688 (.Y(N6768), .A(N6749), .B(N6759));
NAND2BXL inst_cellmath__57_0_I1689 (.Y(N6695), .AN(N6759), .B(N6751));
INVXL inst_cellmath__57_0_I1690 (.Y(N6732), .A(N6768));
NAND4BX1 inst_cellmath__57_0_I1691 (.Y(N6703), .AN(N6767), .B(inst_cellmath__50[19]), .C(inst_cellmath__50[20]), .D(N6768));
NOR2BX1 inst_cellmath__57_0_I1692 (.Y(N6713), .AN(N6731), .B(N6719));
INVXL inst_cellmath__57_0_I1693 (.Y(N6744), .A(N6759));
NOR2XL inst_cellmath__57_0_I1694 (.Y(N6718), .A(N6709), .B(N6759));
INVXL inst_cellmath__57_0_I1695 (.Y(N6762), .A(N6695));
NOR2XL inst_cellmath__57_0_I1696 (.Y(N6758), .A(N6727), .B(N6695));
INVXL inst_cellmath__57_0_I1697 (.Y(N6702), .A(N6732));
NOR2XL inst_cellmath__57_0_I1698 (.Y(N6766), .A(N6767), .B(N6732));
INVXL inst_cellmath__57_0_I1699 (.Y(N6721), .A(N6703));
NAND2XL inst_cellmath__57_0_I1700 (.Y(N6775), .A(inst_cellmath__50[22]), .B(inst_cellmath__50[21]));
NOR2X1 inst_cellmath__57_0_I1701 (.Y(N6777), .A(N6703), .B(N6775));
NOR2BX1 inst_cellmath__57_0_I1702 (.Y(N6701), .AN(inst_cellmath__50[3]), .B(N6776));
NAND2XL inst_cellmath__57_0_I1703 (.Y(N6710), .A(inst_cellmath__50[5]), .B(N6731));
NAND2XL inst_cellmath__57_0_I1704 (.Y(N6748), .A(inst_cellmath__50[7]), .B(N6713));
NAND2XL inst_cellmath__57_0_I1705 (.Y(N6754), .A(inst_cellmath__50[9]), .B(N6744));
NAND2XL inst_cellmath__57_0_I1706 (.Y(N6763), .A(inst_cellmath__50[11]), .B(N6718));
NAND2XL inst_cellmath__57_0_I1707 (.Y(N6729), .A(inst_cellmath__50[13]), .B(N6762));
NAND2XL inst_cellmath__57_0_I1708 (.Y(N6770), .A(inst_cellmath__50[15]), .B(N6758));
NAND2XL inst_cellmath__57_0_I1709 (.Y(N6696), .A(inst_cellmath__50[17]), .B(N6702));
NAND2XL inst_cellmath__57_0_I1710 (.Y(N6705), .A(inst_cellmath__50[19]), .B(N6766));
NAND2XL inst_cellmath__57_0_I1711 (.Y(N6714), .A(inst_cellmath__50[21]), .B(N6721));
NAND2XL inst_cellmath__57_0_I1712 (.Y(N6720), .A(inst_cellmath__50[23]), .B(N6777));
AND3XL inst_cellmath__57_0_I1713 (.Y(inst_cellmath__57[23]), .A(inst_cellmath__50[24]), .B(inst_cellmath__50[23]), .C(N6777));
XOR2XL inst_cellmath__57_0_I1714 (.Y(inst_cellmath__57[0]), .A(inst_cellmath__50[2]), .B(inst_cellmath__55));
XNOR2X1 inst_cellmath__57_0_I1715 (.Y(inst_cellmath__57[1]), .A(N6776), .B(inst_cellmath__50[3]));
XOR2XL inst_cellmath__57_0_I1716 (.Y(inst_cellmath__57[2]), .A(N6701), .B(inst_cellmath__50[4]));
XOR2XL inst_cellmath__57_0_I1717 (.Y(inst_cellmath__57[3]), .A(N6731), .B(inst_cellmath__50[5]));
XNOR2X1 inst_cellmath__57_0_I1718 (.Y(inst_cellmath__57[4]), .A(N6710), .B(inst_cellmath__50[6]));
XOR2XL inst_cellmath__57_0_I1719 (.Y(inst_cellmath__57[5]), .A(N6713), .B(inst_cellmath__50[7]));
XNOR2X1 inst_cellmath__57_0_I1720 (.Y(inst_cellmath__57[6]), .A(N6748), .B(inst_cellmath__50[8]));
XOR2XL inst_cellmath__57_0_I1721 (.Y(inst_cellmath__57[7]), .A(N6744), .B(inst_cellmath__50[9]));
XNOR2X1 inst_cellmath__57_0_I1722 (.Y(inst_cellmath__57[8]), .A(N6754), .B(inst_cellmath__50[10]));
XOR2XL inst_cellmath__57_0_I1723 (.Y(inst_cellmath__57[9]), .A(N6718), .B(inst_cellmath__50[11]));
XNOR2X1 inst_cellmath__57_0_I1724 (.Y(inst_cellmath__57[10]), .A(N6763), .B(inst_cellmath__50[12]));
XOR2XL inst_cellmath__57_0_I1725 (.Y(inst_cellmath__57[11]), .A(N6762), .B(inst_cellmath__50[13]));
XNOR2X1 inst_cellmath__57_0_I1726 (.Y(inst_cellmath__57[12]), .A(N6729), .B(inst_cellmath__50[14]));
XOR2XL inst_cellmath__57_0_I1727 (.Y(inst_cellmath__57[13]), .A(N6758), .B(inst_cellmath__50[15]));
XNOR2X1 inst_cellmath__57_0_I1728 (.Y(inst_cellmath__57[14]), .A(N6770), .B(inst_cellmath__50[16]));
XOR2XL inst_cellmath__57_0_I1729 (.Y(inst_cellmath__57[15]), .A(N6702), .B(inst_cellmath__50[17]));
XNOR2X1 inst_cellmath__57_0_I1730 (.Y(inst_cellmath__57[16]), .A(N6696), .B(inst_cellmath__50[18]));
XOR2XL inst_cellmath__57_0_I1731 (.Y(inst_cellmath__57[17]), .A(N6766), .B(inst_cellmath__50[19]));
XNOR2X1 inst_cellmath__57_0_I1732 (.Y(inst_cellmath__57[18]), .A(N6705), .B(inst_cellmath__50[20]));
XOR2XL inst_cellmath__57_0_I1733 (.Y(inst_cellmath__57[19]), .A(N6721), .B(inst_cellmath__50[21]));
XNOR2X1 inst_cellmath__57_0_I1734 (.Y(inst_cellmath__57[20]), .A(N6714), .B(inst_cellmath__50[22]));
XOR2XL inst_cellmath__57_0_I1735 (.Y(inst_cellmath__57[21]), .A(N6777), .B(inst_cellmath__50[23]));
XNOR2X1 inst_cellmath__57_0_I1736 (.Y(inst_cellmath__57[22]), .A(N6720), .B(inst_cellmath__50[24]));
AOI21XL cynw_cm_float_add2_ieee_I3231 (.Y(N642), .A0(inst_cellmath__45[24]), .A1(inst_cellmath__57[23]), .B0(inst_cellmath__45[25]));
INVXL cynw_cm_float_add2_ieee_I76 (.Y(N574), .A(inst_cellmath__28[8]));
MX2XL inst_cellmath__29_0_I1739 (.Y(inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(N574));
MX2XL inst_cellmath__29_0_I1740 (.Y(inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(N574));
MX2XL inst_cellmath__29_0_I1741 (.Y(inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(N574));
MX2XL inst_cellmath__29_0_I1742 (.Y(inst_cellmath__29[3]), .A(a_exp[3]), .B(N2691), .S0(N574));
MX2XL inst_cellmath__29_0_I1743 (.Y(inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(N574));
MX2XL inst_cellmath__29_0_I1744 (.Y(inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(N574));
MX2XL inst_cellmath__29_0_I1745 (.Y(inst_cellmath__29[6]), .A(a_exp[6]), .B(b_exp[6]), .S0(N574));
MX2XL inst_cellmath__29_0_I1746 (.Y(inst_cellmath__29[7]), .A(a_exp[7]), .B(b_exp[7]), .S0(N574));
NAND3XL inst_cellmath__62_0_I1748 (.Y(N6893), .A(inst_cellmath__29[6]), .B(inst_cellmath__29[7]), .C(inst_cellmath__29[5]));
NOR2XL inst_cellmath__62_0_I1749 (.Y(N6892), .A(inst_cellmath__29[0]), .B(N6893));
NAND3XL inst_cellmath__62_0_I1750 (.Y(N6889), .A(inst_cellmath__29[4]), .B(inst_cellmath__29[3]), .C(N6892));
NAND3BXL inst_cellmath__62_0_I3232 (.Y(N6883), .AN(N6889), .B(inst_cellmath__29[1]), .C(inst_cellmath__29[2]));
NOR2XL inst_cellmath__62_0_I1752 (.Y(inst_cellmath__62), .A(N6883), .B(N642));
ADDHX1 inst_cellmath__59_0_I1756 (.CO(N6931), .S(N6918), .A(inst_cellmath__29[1]), .B(inst_cellmath__29[2]));
ADDHX1 inst_cellmath__59_0_I1757 (.CO(N6902), .S(N6944), .A(inst_cellmath__29[3]), .B(N6931));
ADDHX1 inst_cellmath__59_0_I1758 (.CO(N6923), .S(N6911), .A(inst_cellmath__29[4]), .B(N6902));
INVXL inst_cellmath__59_0_I1759 (.Y(N6936), .A(inst_cellmath__29[5]));
INVXL inst_cellmath__59_0_I1760 (.Y(N6928), .A(inst_cellmath__29[6]));
INVXL inst_cellmath__59_0_I1761 (.Y(N6921), .A(inst_cellmath__29[7]));
NOR2XL inst_cellmath__59_0_I1762 (.Y(N6941), .A(inst_cellmath__29[0]), .B(inst_cellmath__57[23]));
CLKXOR2X1 inst_cellmath__59_0_I3234 (.Y(N6951), .A(inst_cellmath__29[0]), .B(inst_cellmath__57[23]));
NAND2XL inst_cellmath__59_0_I1764 (.Y(N6909), .A(inst_cellmath__29[1]), .B(inst_cellmath__49[1]));
XNOR2X1 inst_cellmath__59_0_I1765 (.Y(N6919), .A(inst_cellmath__29[1]), .B(inst_cellmath__49[1]));
XOR2XL inst_cellmath__59_0_I1766 (.Y(N6946), .A(N6918), .B(N6360));
XNOR2X1 inst_cellmath__59_0_I1767 (.Y(N6913), .A(N6944), .B(N6439));
XOR2XL inst_cellmath__59_0_I1768 (.Y(N6938), .A(N6911), .B(N6311));
XNOR2X1 inst_cellmath__59_0_I1769 (.Y(N6908), .A(N6936), .B(N6923));
XOR2XL inst_cellmath__59_0_I1770 (.Y(N6929), .A(inst_cellmath__29[5]), .B(N6928));
XNOR2X1 inst_cellmath__59_0_I1771 (.Y(N6901), .A(inst_cellmath__29[6]), .B(N6921));
AOI21X1 inst_cellmath__59_0_I1772 (.Y(N6948), .A0(inst_cellmath__49[0]), .A1(N6951), .B0(N6941));
OAI21X1 inst_cellmath__59_0_I1773 (.Y(N6933), .A0(N6919), .A1(N6948), .B0(N6909));
AOI2BB2X2 inst_cellmath__59_0_I1774 (.Y(N6917), .A0N(N6918), .A1N(N6360), .B0(N6933), .B1(N6946));
OAI22X2 inst_cellmath__59_0_I1775 (.Y(N6954), .A0(N6913), .A1(N6917), .B0(N6944), .B1(N6439));
AOI2BB2X2 inst_cellmath__59_0_I1776 (.Y(N6932), .A0N(N6911), .A1N(N6311), .B0(N6954), .B1(N6938));
OAI22X2 inst_cellmath__59_0_I1777 (.Y(N6905), .A0(N6908), .A1(N6932), .B0(N6936), .B1(N6923));
AOI2BB2X2 inst_cellmath__59_0_I1778 (.Y(N6930), .A0N(inst_cellmath__29[5]), .A1N(N6928), .B0(N6905), .B1(N6929));
OAI22X2 inst_cellmath__59_0_I1779 (.Y(N6950), .A0(N6901), .A1(N6930), .B0(inst_cellmath__29[6]), .B1(N6921));
XNOR2X1 inst_cellmath__59_0_I3092 (.Y(N8785), .A(inst_cellmath__49[0]), .B(N6951));
XNOR2X1 inst_cellmath__59_0_I1781 (.Y(inst_cellmath__59[1]), .A(N6948), .B(N6919));
XNOR2X1 inst_cellmath__59_0_I1782 (.Y(inst_cellmath__59[2]), .A(N6933), .B(N6946));
XNOR2X1 inst_cellmath__59_0_I1783 (.Y(inst_cellmath__59[3]), .A(N6917), .B(N6913));
XNOR2X1 inst_cellmath__59_0_I1784 (.Y(inst_cellmath__59[4]), .A(N6954), .B(N6938));
XNOR2X1 inst_cellmath__59_0_I1785 (.Y(inst_cellmath__59[5]), .A(N6932), .B(N6908));
XNOR2X1 inst_cellmath__59_0_I1786 (.Y(inst_cellmath__59[6]), .A(N6905), .B(N6929));
XNOR2X1 inst_cellmath__59_0_I1787 (.Y(inst_cellmath__59[7]), .A(N6930), .B(N6901));
XNOR2X1 inst_cellmath__59_0_I1788 (.Y(inst_cellmath__59[8]), .A(N6950), .B(N6921));
AND2XL inst_cellmath__59_0_I1789 (.Y(inst_cellmath__59[9]), .A(N6921), .B(N6950));
NOR3XL inst_cellmath__60__44__I1791 (.Y(N6999), .A(N8785), .B(inst_cellmath__59[1]), .C(inst_cellmath__59[3]));
NOR2XL inst_cellmath__60__44__I1793 (.Y(N6997), .A(inst_cellmath__59[7]), .B(inst_cellmath__59[8]));
NAND2XL inst_cellmath__60__44__I1794 (.Y(N7000), .A(N6997), .B(N6999));
OR4X1 inst_cellmath__60__44__I7946 (.Y(N8722), .A(inst_cellmath__59[2]), .B(inst_cellmath__59[4]), .C(inst_cellmath__59[5]), .D(inst_cellmath__59[6]));
OR4X1 inst_cellmath__71_1_I1796 (.Y(N7018), .A(N706), .B(inst_cellmath__12), .C(inst_cellmath__17), .D(inst_cellmath__63));
NOR4X1 inst_cellmath__71_1_I1797 (.Y(N7020), .A(N7018), .B(inst_cellmath__49[5]), .C(inst_cellmath__62), .D(inst_cellmath__59[9]));
OR4X1 cynw_cm_float_add2_ieee_I3238 (.Y(N650), .A(inst_cellmath__4), .B(inst_cellmath__8), .C(N635), .D(N634));
AND2XL cynw_cm_float_add2_ieee_I1802 (.Y(N651), .A(N650), .B(inst_cellmath__62));
OR4X1 cynw_cm_float_add2_ieee_I1803 (.Y(inst_cellmath__68[0]), .A(inst_cellmath__12), .B(inst_cellmath__17), .C(inst_cellmath__63), .D(N651));
OR4X1 inst_cellmath__72_0_I3239 (.Y(N7068), .A(inst_cellmath__12), .B(inst_cellmath__17), .C(inst_cellmath__63), .D(inst_cellmath__62));
OA21X1 inst_cellmath__72_0_I3240 (.Y(N7074), .A0(N8722), .A1(N7000), .B0(N7020));
INVXL inst_cellmath__72_0_I1808 (.Y(N7056), .A(N7074));
MX2XL inst_cellmath__72_0_I1809 (.Y(x[23]), .A(N8785), .B(inst_cellmath__68[0]), .S0(N7056));
MX2XL inst_cellmath__72_0_I1810 (.Y(x[24]), .A(inst_cellmath__59[1]), .B(N7068), .S0(N7056));
MX2XL inst_cellmath__72_0_I1811 (.Y(x[25]), .A(inst_cellmath__59[2]), .B(N7068), .S0(N7056));
MX2XL inst_cellmath__72_0_I1812 (.Y(x[26]), .A(inst_cellmath__59[3]), .B(N7068), .S0(N7056));
MX2XL inst_cellmath__72_0_I1813 (.Y(x[27]), .A(inst_cellmath__59[4]), .B(N7068), .S0(N7056));
MX2XL inst_cellmath__72_0_I1814 (.Y(x[28]), .A(inst_cellmath__59[5]), .B(N7068), .S0(N7056));
MX2XL inst_cellmath__72_0_I1815 (.Y(x[29]), .A(inst_cellmath__59[6]), .B(N7068), .S0(N7056));
MX2XL inst_cellmath__72_0_I1816 (.Y(x[30]), .A(inst_cellmath__59[7]), .B(N7068), .S0(N7056));
NAND2XL inst_cellmath__7_0_I1817 (.Y(N7092), .A(rm[0]), .B(rm[1]));
NOR2XL inst_cellmath__7_0_I1818 (.Y(inst_cellmath__7), .A(rm[2]), .B(N7092));
XNOR2X1 cynw_cm_float_add2_ieee_I1819 (.Y(N652), .A(inst_cellmath__48), .B(inst_cellmath__5));
OR2XL cynw_cm_float_add2_ieee_I1820 (.Y(N653), .A(inst_cellmath__7), .B(N652));
NOR3BXL inst_cellmath__70_0_I1821 (.Y(N7111), .AN(N653), .B(inst_cellmath__8), .C(inst_cellmath__4));
AND2XL inst_cellmath__70_0_I1822 (.Y(inst_cellmath__70), .A(N7111), .B(inst_cellmath__62));
INVX2 inst_cellmath__73_0_I3190 (.Y(N8825), .A(N7074));
INVX3 inst_cellmath__73_0_I3195 (.Y(N8830), .A(N8825));
INVX1 inst_cellmath__73_0_I7908 (.Y(N13892), .A(N8830));
INVX3 inst_cellmath__73_0_I7909 (.Y(N13893), .A(N13892));
INVXL inst_cellmath__73_0_I3191 (.Y(N8826), .A(N8825));
NOR2X8 inst_cellmath__73_0_I1824 (.Y(N7150), .A(inst_cellmath__63), .B(N8830));
NOR2BX2 inst_cellmath__73_0_I1825 (.Y(N7141), .AN(inst_cellmath__63), .B(N7074));
AOI22XL inst_cellmath__73_0_I1826 (.Y(N7125), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[0]));
AOI22XL inst_cellmath__73_0_I1827 (.Y(N7169), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[1]));
AOI22XL inst_cellmath__73_0_I1828 (.Y(N7210), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[2]));
AOI22XL inst_cellmath__73_0_I1829 (.Y(N7156), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[3]));
AOI22XL inst_cellmath__73_0_I1830 (.Y(N7198), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[4]));
AOI22XL inst_cellmath__73_0_I1831 (.Y(N7142), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[5]));
AOI22XL inst_cellmath__73_0_I1832 (.Y(N7186), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[6]));
AOI22XL inst_cellmath__73_0_I1833 (.Y(N7129), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[7]));
AOI22XL inst_cellmath__73_0_I1834 (.Y(N7173), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[8]));
AOI22XL inst_cellmath__73_0_I1835 (.Y(N7117), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[9]));
AOI22XL inst_cellmath__73_0_I1836 (.Y(N7161), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[10]));
AOI22XL inst_cellmath__73_0_I1837 (.Y(N7202), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[11]));
AOI22XL inst_cellmath__73_0_I1838 (.Y(N7146), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[12]));
AOI22XL inst_cellmath__73_0_I1839 (.Y(N7190), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[13]));
AOI22XL inst_cellmath__73_0_I1840 (.Y(N7133), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[14]));
AOI22X1 inst_cellmath__73_0_I1841 (.Y(N7178), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[15]));
AOI22XL inst_cellmath__73_0_I1842 (.Y(N7122), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[16]));
AOI22XL inst_cellmath__73_0_I1843 (.Y(N7166), .A0(inst_cellmath__70), .A1(N7150), .B0(N13893), .B1(inst_cellmath__57[17]));
AOI22XL inst_cellmath__73_0_I1844 (.Y(N7207), .A0(inst_cellmath__70), .A1(N7150), .B0(N8826), .B1(inst_cellmath__57[18]));
AOI22XL inst_cellmath__73_0_I1845 (.Y(N7153), .A0(inst_cellmath__70), .A1(N7150), .B0(N8826), .B1(inst_cellmath__57[19]));
AOI22XL inst_cellmath__73_0_I1846 (.Y(N7195), .A0(inst_cellmath__70), .A1(N7150), .B0(N8826), .B1(inst_cellmath__57[20]));
AOI22XL inst_cellmath__73_0_I1847 (.Y(N7138), .A0(inst_cellmath__70), .A1(N7150), .B0(N8826), .B1(inst_cellmath__57[21]));
AOI22XL inst_cellmath__73_0_I1848 (.Y(N7182), .A0(inst_cellmath__70), .A1(N7150), .B0(N8826), .B1(inst_cellmath__57[22]));
OAI2BB1XL inst_cellmath__73_0_I1849 (.Y(x[0]), .A0N(N7141), .A1N(inst_cellmath__64[0]), .B0(N7125));
OAI2BB1XL inst_cellmath__73_0_I1850 (.Y(x[1]), .A0N(N7141), .A1N(inst_cellmath__64[1]), .B0(N7169));
OAI2BB1XL inst_cellmath__73_0_I1851 (.Y(x[2]), .A0N(N7141), .A1N(inst_cellmath__64[2]), .B0(N7210));
OAI2BB1XL inst_cellmath__73_0_I1852 (.Y(x[3]), .A0N(N7141), .A1N(inst_cellmath__64[3]), .B0(N7156));
OAI2BB1XL inst_cellmath__73_0_I1853 (.Y(x[4]), .A0N(N7141), .A1N(inst_cellmath__64[4]), .B0(N7198));
OAI2BB1XL inst_cellmath__73_0_I1854 (.Y(x[5]), .A0N(N7141), .A1N(inst_cellmath__64[5]), .B0(N7142));
OAI2BB1XL inst_cellmath__73_0_I1855 (.Y(x[6]), .A0N(N7141), .A1N(inst_cellmath__64[6]), .B0(N7186));
OAI2BB1XL inst_cellmath__73_0_I1856 (.Y(x[7]), .A0N(N7141), .A1N(inst_cellmath__64[7]), .B0(N7129));
OAI2BB1XL inst_cellmath__73_0_I1857 (.Y(x[8]), .A0N(N7141), .A1N(inst_cellmath__64[8]), .B0(N7173));
OAI2BB1XL inst_cellmath__73_0_I1858 (.Y(x[9]), .A0N(N7141), .A1N(inst_cellmath__64[9]), .B0(N7117));
OAI2BB1XL inst_cellmath__73_0_I1859 (.Y(x[10]), .A0N(N7141), .A1N(inst_cellmath__64[10]), .B0(N7161));
OAI2BB1XL inst_cellmath__73_0_I1860 (.Y(x[11]), .A0N(N7141), .A1N(inst_cellmath__64[11]), .B0(N7202));
OAI2BB1XL inst_cellmath__73_0_I1861 (.Y(x[12]), .A0N(N7141), .A1N(inst_cellmath__64[12]), .B0(N7146));
OAI2BB1XL inst_cellmath__73_0_I1862 (.Y(x[13]), .A0N(N7141), .A1N(inst_cellmath__64[13]), .B0(N7190));
OAI2BB1XL inst_cellmath__73_0_I1863 (.Y(x[14]), .A0N(N7141), .A1N(inst_cellmath__64[14]), .B0(N7133));
OAI2BB1X1 inst_cellmath__73_0_I1864 (.Y(x[15]), .A0N(N7141), .A1N(inst_cellmath__64[15]), .B0(N7178));
OAI2BB1XL inst_cellmath__73_0_I1865 (.Y(x[16]), .A0N(N7141), .A1N(inst_cellmath__64[16]), .B0(N7122));
OAI2BB1XL inst_cellmath__73_0_I1866 (.Y(x[17]), .A0N(N7141), .A1N(inst_cellmath__64[17]), .B0(N7166));
OAI2BB1XL inst_cellmath__73_0_I1867 (.Y(x[18]), .A0N(N7141), .A1N(inst_cellmath__64[18]), .B0(N7207));
OAI2BB1XL inst_cellmath__73_0_I1868 (.Y(x[19]), .A0N(N7141), .A1N(inst_cellmath__64[19]), .B0(N7153));
OAI2BB1XL inst_cellmath__73_0_I1869 (.Y(x[20]), .A0N(N7141), .A1N(inst_cellmath__64[20]), .B0(N7195));
OAI2BB1XL inst_cellmath__73_0_I1870 (.Y(x[21]), .A0N(N7141), .A1N(inst_cellmath__64[21]), .B0(N7138));
NAND2BXL inst_cellmath__73_0_I1871 (.Y(x[22]), .AN(N7141), .B(N7182));
assign inst_cellmath__28[0] = 1'B0;
assign inst_cellmath__28[1] = 1'B0;
assign inst_cellmath__28[2] = 1'B0;
assign inst_cellmath__28[3] = 1'B0;
assign inst_cellmath__28[4] = 1'B0;
assign inst_cellmath__28[5] = 1'B0;
assign inst_cellmath__28[6] = 1'B0;
assign inst_cellmath__28[7] = 1'B0;
assign inst_cellmath__33[0] = 1'B0;
assign inst_cellmath__33[1] = 1'B0;
assign inst_cellmath__33[2] = 1'B0;
assign inst_cellmath__33[3] = 1'B0;
assign inst_cellmath__33[4] = 1'B0;
assign inst_cellmath__33[5] = 1'B0;
assign inst_cellmath__33[6] = 1'B0;
assign inst_cellmath__33[7] = 1'B0;
assign inst_cellmath__33[8] = 1'B0;
assign inst_cellmath__33[9] = 1'B0;
assign inst_cellmath__33[10] = 1'B0;
assign inst_cellmath__33[11] = 1'B0;
assign inst_cellmath__33[12] = 1'B0;
assign inst_cellmath__33[13] = 1'B0;
assign inst_cellmath__33[14] = 1'B0;
assign inst_cellmath__33[15] = 1'B0;
assign inst_cellmath__33[16] = 1'B0;
assign inst_cellmath__33[17] = 1'B0;
assign inst_cellmath__33[18] = 1'B0;
assign inst_cellmath__33[19] = 1'B0;
assign inst_cellmath__33[20] = 1'B0;
assign inst_cellmath__33[21] = 1'B0;
assign inst_cellmath__33[22] = 1'B0;
assign inst_cellmath__33[23] = 1'B0;
assign inst_cellmath__33[26] = 1'B0;
assign inst_cellmath__33[28] = 1'B0;
assign inst_cellmath__33[32] = 1'B0;
assign inst_cellmath__33[34] = 1'B0;
assign inst_cellmath__35[1] = 1'B0;
assign inst_cellmath__36[0] = 1'B0;
assign inst_cellmath__36[1] = 1'B0;
assign inst_cellmath__36[2] = 1'B0;
assign inst_cellmath__36[3] = 1'B0;
assign inst_cellmath__36[4] = 1'B0;
assign inst_cellmath__36[5] = 1'B0;
assign inst_cellmath__36[6] = 1'B0;
assign inst_cellmath__36[7] = 1'B0;
assign inst_cellmath__36[8] = 1'B0;
assign inst_cellmath__36[9] = 1'B0;
assign inst_cellmath__36[10] = 1'B0;
assign inst_cellmath__36[11] = 1'B0;
assign inst_cellmath__36[12] = 1'B0;
assign inst_cellmath__36[13] = 1'B0;
assign inst_cellmath__36[14] = 1'B0;
assign inst_cellmath__36[15] = 1'B0;
assign inst_cellmath__36[16] = 1'B0;
assign inst_cellmath__36[17] = 1'B0;
assign inst_cellmath__36[18] = 1'B0;
assign inst_cellmath__36[19] = 1'B0;
assign inst_cellmath__36[20] = 1'B0;
assign inst_cellmath__36[21] = 1'B0;
assign inst_cellmath__36[22] = 1'B0;
assign inst_cellmath__36[23] = 1'B0;
assign inst_cellmath__36[24] = 1'B0;
assign inst_cellmath__36[25] = 1'B0;
assign inst_cellmath__36[49] = 1'B1;
assign inst_cellmath__37[42] = 1'B0;
assign inst_cellmath__37[43] = 1'B0;
assign inst_cellmath__37[44] = 1'B0;
assign inst_cellmath__37[45] = 1'B0;
assign inst_cellmath__37[46] = 1'B0;
assign inst_cellmath__37[47] = 1'B0;
assign inst_cellmath__37[48] = 1'B0;
assign inst_cellmath__45[26] = 1'B0;
assign inst_cellmath__49[2] = 1'B0;
assign inst_cellmath__49[3] = 1'B0;
assign inst_cellmath__49[4] = 1'B0;
assign inst_cellmath__50[0] = 1'B0;
assign inst_cellmath__59[0] = 1'B0;
assign inst_cellmath__64[22] = 1'B1;
assign inst_cellmath__68[1] = 1'B0;
assign inst_cellmath__68[2] = 1'B0;
assign inst_cellmath__68[3] = 1'B0;
assign inst_cellmath__68[4] = 1'B0;
assign inst_cellmath__68[5] = 1'B0;
assign inst_cellmath__68[6] = 1'B0;
assign inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  urPwSAjbqx4= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



