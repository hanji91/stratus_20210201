/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:25:22 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_5 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895;
wire N5527,N5534,N5541,N5548,N5555,N5562,N5569 
	,N5576,N5583,N5590,N5597,N5604,N5611,N5618,N5625 
	,N5632,N5639,N5646,N5653,N5660,N5667,N5679,N5738 
	,N5740,N5976,N5989,N5991,N6015,N6017,N6024,N6031 
	,N6038,N6045,N6052,N6059,N6066,N6073,N6080,N6087 
	,N6094,N6101,N6108,N6115,N6122,N6129,N6136,N6143 
	,N6157,N6176,N6183,N6190,N6197,N6199,N6206,N6213 
	,N6220,N6227,N6311,N6316,N6436,N6442,N6451,N6460 
	,N6469,N6478,N6487,N6496,N6505,N6514,N6523,N6532 
	,N6541,N6550,N6559,N6568,N6577,N6586,N6595,N6604 
	,N6613,N6622,N6631,N6640,N6667,N6875,N6915,N6921 
	,N6946,N6959,N6962,N6964,N6966,N6982,N6988,N7029 
	,N7035,N7044,N7050,N7058,N7060,N7066,N7076,N7078 
	,N7088,N7096,N7114,N7148,N7159,N7908,N7910,N7912 
	,N7934,N8072,N8357,N8377,N8595,N8597,N8599,N9114 
	,N9122,N9129,N9144,N9151,N9158,N9166,N9173,N9180 
	,N9187,N9195,N9203,N9211,N9219,N9227,N9235,N9243 
	,N9251,N9259,N9267,N9273,N9275,N9281,N9283,N9289 
	,N9291,N9294,N9301,N9313,N9320,N9327,N9329,N9334 
	,N9336,N9341,N9348,N9355,N9357,N9362,N9370,N9372 
	,N9374,N9380,N9388,N9390,N9396,N9398,N9416,N9418 
	,N9437,N9439,N9457,N9459,N9467,N9469,N9489,N9493 
	,N9497,N9501,N9982,N9985,N9988,N10010,N10012,N10015 
	,N10416,N10417,N10418,N10419;
reg x_reg_L0_15__retimed_I5178_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5178_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664;
	end
assign N10015 = x_reg_L0_15__retimed_I5178_QOUT;
reg x_reg_L0_15__retimed_I5177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5177_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814;
	end
assign N10012 = x_reg_L0_15__retimed_I5177_QOUT;
reg x_reg_L0_15__retimed_I5176_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5176_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725;
	end
assign N10010 = x_reg_L0_15__retimed_I5176_QOUT;
reg x_reg_L0_15__retimed_I5167_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5167_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839;
	end
assign N9988 = x_reg_L0_15__retimed_I5167_QOUT;
reg x_reg_L0_15__retimed_I5166_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5166_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686;
	end
assign N9985 = x_reg_L0_15__retimed_I5166_QOUT;
reg x_reg_L0_15__retimed_I5165_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5165_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816;
	end
assign N9982 = x_reg_L0_15__retimed_I5165_QOUT;
reg x_reg_L1_17__retimed_I4959_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4959_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5];
	end
assign N9501 = x_reg_L1_17__retimed_I4959_QOUT;
reg x_reg_L1_17__retimed_I4957_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4957_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930;
	end
assign N9497 = x_reg_L1_17__retimed_I4957_QOUT;
reg x_reg_L1_17__retimed_I4955_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4955_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4];
	end
assign N9493 = x_reg_L1_17__retimed_I4955_QOUT;
reg x_reg_L1_17__retimed_I4953_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4953_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905;
	end
assign N9489 = x_reg_L1_17__retimed_I4953_QOUT;
reg x_reg_L0_15__retimed_I4943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4943_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771;
	end
assign N9469 = x_reg_L0_15__retimed_I4943_QOUT;
reg x_reg_L0_15__retimed_I4942_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4942_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728;
	end
assign N9467 = x_reg_L0_15__retimed_I4942_QOUT;
reg x_reg_L0_15__retimed_I4940_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4940_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698;
	end
assign N9459 = x_reg_L0_15__retimed_I4940_QOUT;
reg x_reg_L0_15__retimed_I4939_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4939_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655;
	end
assign N9457 = x_reg_L0_15__retimed_I4939_QOUT;
reg x_reg_L0_15__retimed_I4933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4933_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836;
	end
assign N9439 = x_reg_L0_15__retimed_I4933_QOUT;
reg x_reg_L0_15__retimed_I4932_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4932_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790;
	end
assign N9437 = x_reg_L0_15__retimed_I4932_QOUT;
reg x_reg_L0_15__retimed_I4926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4926_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660;
	end
assign N9418 = x_reg_L0_15__retimed_I4926_QOUT;
reg x_reg_L0_15__retimed_I4925_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4925_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813;
	end
assign N9416 = x_reg_L0_15__retimed_I4925_QOUT;
reg x_reg_L0_15__retimed_I4920_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4920_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805;
	end
assign N9398 = x_reg_L0_15__retimed_I4920_QOUT;
reg x_reg_L0_15__retimed_I4919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4919_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759;
	end
assign N9396 = x_reg_L0_15__retimed_I4919_QOUT;
reg x_reg_L0_15__retimed_I4917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4917_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811;
	end
assign N9390 = x_reg_L0_15__retimed_I4917_QOUT;
reg x_reg_L0_15__retimed_I4916_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4916_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659;
	end
assign N9388 = x_reg_L0_15__retimed_I4916_QOUT;
reg x_reg_L0_15__retimed_I4913_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4913_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734;
	end
assign N9380 = x_reg_L0_15__retimed_I4913_QOUT;
reg x_reg_L0_15__retimed_I4911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4911_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778;
	end
assign N9374 = x_reg_L0_15__retimed_I4911_QOUT;
reg x_reg_L0_15__retimed_I4910_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4910_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671;
	end
assign N9372 = x_reg_L0_15__retimed_I4910_QOUT;
reg x_reg_L0_15__retimed_I4909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4909_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777;
	end
assign N9370 = x_reg_L0_15__retimed_I4909_QOUT;
reg x_reg_L0_15__retimed_I4906_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4906_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832;
	end
assign N9362 = x_reg_L0_15__retimed_I4906_QOUT;
reg x_reg_L0_15__retimed_I4904_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4904_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744;
	end
assign N9357 = x_reg_L0_15__retimed_I4904_QOUT;
reg x_reg_L0_15__retimed_I4903_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4903_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788;
	end
assign N9355 = x_reg_L0_15__retimed_I4903_QOUT;
reg x_reg_L0_15__retimed_I4900_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4900_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779;
	end
assign N9348 = x_reg_L0_15__retimed_I4900_QOUT;
reg x_reg_L0_15__retimed_I4897_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4897_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753;
	end
assign N9341 = x_reg_L0_15__retimed_I4897_QOUT;
reg x_reg_L0_15__retimed_I4895_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4895_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756;
	end
assign N9336 = x_reg_L0_15__retimed_I4895_QOUT;
reg x_reg_L0_15__retimed_I4894_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4894_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800;
	end
assign N9334 = x_reg_L0_15__retimed_I4894_QOUT;
reg x_reg_L0_15__retimed_I4892_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4892_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819;
	end
assign N9329 = x_reg_L0_15__retimed_I4892_QOUT;
reg x_reg_L0_15__retimed_I4891_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4891_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666;
	end
assign N9327 = x_reg_L0_15__retimed_I4891_QOUT;
reg x_reg_L0_15__retimed_I4888_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4888_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682;
	end
assign N9320 = x_reg_L0_15__retimed_I4888_QOUT;
reg x_reg_L0_15__retimed_I4885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4885_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829;
	end
assign N9313 = x_reg_L0_15__retimed_I4885_QOUT;
reg x_reg_L0_15__retimed_I4880_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4880_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656;
	end
assign N9301 = x_reg_L0_15__retimed_I4880_QOUT;
reg x_reg_L0_15__retimed_I4877_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4877_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801;
	end
assign N9294 = x_reg_L0_15__retimed_I4877_QOUT;
reg x_reg_L0_15__retimed_I4876_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4876_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703;
	end
assign N9291 = x_reg_L0_15__retimed_I4876_QOUT;
reg x_reg_L0_15__retimed_I4875_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4875_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668;
	end
assign N9289 = x_reg_L0_15__retimed_I4875_QOUT;
reg x_reg_L0_15__retimed_I4874_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4874_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786;
	end
assign N9283 = x_reg_L0_15__retimed_I4874_QOUT;
reg x_reg_L0_15__retimed_I4873_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4873_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796;
	end
assign N9281 = x_reg_L0_15__retimed_I4873_QOUT;
reg x_reg_L0_15__retimed_I4872_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4872_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680;
	end
assign N9275 = x_reg_L0_15__retimed_I4872_QOUT;
reg x_reg_L0_15__retimed_I4871_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4871_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643;
	end
assign N9273 = x_reg_L0_15__retimed_I4871_QOUT;
reg x_reg_L0_15__retimed_I4870_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4870_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760;
	end
assign N9267 = x_reg_L0_15__retimed_I4870_QOUT;
reg x_reg_L0_15__retimed_I4868_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4868_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652;
	end
assign N9259 = x_reg_L0_15__retimed_I4868_QOUT;
reg x_reg_L0_15__retimed_I4866_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4866_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824;
	end
assign N9251 = x_reg_L0_15__retimed_I4866_QOUT;
reg x_reg_L0_15__retimed_I4864_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4864_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711;
	end
assign N9243 = x_reg_L0_15__retimed_I4864_QOUT;
reg x_reg_L0_15__retimed_I4862_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4862_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735;
	end
assign N9235 = x_reg_L0_15__retimed_I4862_QOUT;
reg x_reg_L0_15__retimed_I4860_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4860_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798;
	end
assign N9227 = x_reg_L0_15__retimed_I4860_QOUT;
reg x_reg_L0_15__retimed_I4858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4858_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772;
	end
assign N9219 = x_reg_L0_15__retimed_I4858_QOUT;
reg x_reg_L0_15__retimed_I4856_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4856_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689;
	end
assign N9211 = x_reg_L0_15__retimed_I4856_QOUT;
reg x_reg_L0_15__retimed_I4854_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4854_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
	end
assign N9203 = x_reg_L0_15__retimed_I4854_QOUT;
reg x_reg_L0_15__retimed_I4852_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4852_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721;
	end
assign N9195 = x_reg_L0_15__retimed_I4852_QOUT;
reg x_reg_L0_15__retimed_I4850_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4850_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809;
	end
assign N9187 = x_reg_L0_15__retimed_I4850_QOUT;
reg x_reg_L0_15__retimed_I4848_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4848_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675;
	end
assign N9180 = x_reg_L0_15__retimed_I4848_QOUT;
reg x_reg_L0_15__retimed_I4846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4846_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700;
	end
assign N9173 = x_reg_L0_15__retimed_I4846_QOUT;
reg x_reg_L0_15__retimed_I4844_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4844_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665;
	end
assign N9166 = x_reg_L0_15__retimed_I4844_QOUT;
reg x_reg_L0_15__retimed_I4842_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4842_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758;
	end
assign N9158 = x_reg_L0_15__retimed_I4842_QOUT;
reg x_reg_L0_15__retimed_I4840_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4840_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648;
	end
assign N9151 = x_reg_L0_15__retimed_I4840_QOUT;
reg x_reg_L0_15__retimed_I4838_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4838_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24];
	end
assign N9144 = x_reg_L0_15__retimed_I4838_QOUT;
reg x_reg_L0_15__retimed_I4834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4834_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783;
	end
assign N9129 = x_reg_L0_15__retimed_I4834_QOUT;
reg x_reg_L0_15__retimed_I4832_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4832_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837;
	end
assign N9122 = x_reg_L0_15__retimed_I4832_QOUT;
reg x_reg_L0_15__retimed_I4830_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4830_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731;
	end
assign N9114 = x_reg_L0_15__retimed_I4830_QOUT;
reg x_reg_L0_15__retimed_I4668_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4668_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630;
	end
assign N8599 = x_reg_L0_15__retimed_I4668_QOUT;
reg x_reg_L0_15__retimed_I4667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4667_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24];
	end
assign N8597 = x_reg_L0_15__retimed_I4667_QOUT;
reg x_reg_L0_15__retimed_I4666_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4666_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
	end
assign N8595 = x_reg_L0_15__retimed_I4666_QOUT;
reg x_reg_L0_15__retimed_I4614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4614_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N8377 = x_reg_L0_15__retimed_I4614_QOUT;
reg x_reg_L0_15__retimed_I4606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4606_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
	end
assign N8357 = x_reg_L0_15__retimed_I4606_QOUT;
reg x_reg_L0_15__retimed_I4517_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4517_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4;
	end
assign N8072 = x_reg_L0_15__retimed_I4517_QOUT;
reg x_reg_L0_15__retimed_I4468_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4468_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638;
	end
assign N7934 = x_reg_L0_15__retimed_I4468_QOUT;
reg x_reg_L0_15__retimed_I4459_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4459_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
	end
assign N7912 = x_reg_L0_15__retimed_I4459_QOUT;
reg x_reg_L0_15__retimed_I4458_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4458_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635;
	end
assign N7910 = x_reg_L0_15__retimed_I4458_QOUT;
reg x_reg_L0_15__retimed_I4457_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4457_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N7908 = x_reg_L0_15__retimed_I4457_QOUT;
reg x_reg_L0_15__retimed_I4165_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4165_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0];
	end
assign N7159 = x_reg_L0_15__retimed_I4165_QOUT;
reg x_reg_L0_15__retimed_I4161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4161_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
	end
assign N7148 = x_reg_L0_15__retimed_I4161_QOUT;
reg x_reg_L0_15__retimed_I4149_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4149_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918;
	end
assign N7114 = x_reg_L0_15__retimed_I4149_QOUT;
reg x_reg_L0_15__retimed_I4142_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4142_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944;
	end
assign N7096 = x_reg_L0_15__retimed_I4142_QOUT;
reg x_reg_L0_15__retimed_I4139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4139_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911;
	end
assign N7088 = x_reg_L0_15__retimed_I4139_QOUT;
reg x_reg_L0_15__retimed_I4135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4135_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923;
	end
assign N7078 = x_reg_L0_15__retimed_I4135_QOUT;
reg x_reg_L0_15__retimed_I4134_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4134_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936;
	end
assign N7076 = x_reg_L0_15__retimed_I4134_QOUT;
reg x_reg_L1_17__retimed_I4130_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4130_QOUT <= N7035;
	end
assign N7066 = x_reg_L1_17__retimed_I4130_QOUT;
reg x_reg_L0_15__retimed_I4128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4128_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928;
	end
assign N7060 = x_reg_L0_15__retimed_I4128_QOUT;
reg x_reg_L0_15__retimed_I4127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4127_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
	end
assign N7058 = x_reg_L0_15__retimed_I4127_QOUT;
reg x_reg_L1_17__retimed_I4124_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4124_QOUT <= N6988;
	end
assign N7050 = x_reg_L1_17__retimed_I4124_QOUT;
reg x_reg_L1_17__retimed_I4122_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4122_QOUT <= N6982;
	end
assign N7044 = x_reg_L1_17__retimed_I4122_QOUT;
reg x_reg_L0_15__retimed_I4118_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4118_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
	end
assign N7035 = x_reg_L0_15__retimed_I4118_QOUT;
reg x_reg_L1_17__retimed_I4116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4116_QOUT <= N6915;
	end
assign N7029 = x_reg_L1_17__retimed_I4116_QOUT;
reg x_reg_L0_15__retimed_I4101_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4101_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901;
	end
assign N6988 = x_reg_L0_15__retimed_I4101_QOUT;
reg x_reg_L0_15__retimed_I4099_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4099_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921;
	end
assign N6982 = x_reg_L0_15__retimed_I4099_QOUT;
reg x_reg_L1_17__retimed_I4092_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4092_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
	end
assign N6966 = x_reg_L1_17__retimed_I4092_QOUT;
reg x_reg_L1_17__retimed_I4091_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4091_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5];
	end
assign N6964 = x_reg_L1_17__retimed_I4091_QOUT;
reg x_reg_L1_17__retimed_I4090_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4090_QOUT <= N6875;
	end
assign N6962 = x_reg_L1_17__retimed_I4090_QOUT;
reg x_reg_L1_17__retimed_I4089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I4089_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999;
	end
assign N6959 = x_reg_L1_17__retimed_I4089_QOUT;
reg x_reg_L0_15__retimed_I4084_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4084_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883;
	end
assign N6946 = x_reg_L0_15__retimed_I4084_QOUT;
reg x_reg_L0_15__retimed_I4076_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4076_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908;
	end
assign N6921 = x_reg_L0_15__retimed_I4076_QOUT;
reg x_reg_L0_15__retimed_I4074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4074_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929;
	end
assign N6915 = x_reg_L0_15__retimed_I4074_QOUT;
reg x_reg_L0_15__retimed_I4058_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I4058_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018;
	end
assign N6875 = x_reg_L0_15__retimed_I4058_QOUT;
reg x_reg_L1_22__retimed_I4004_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I4004_QOUT <= N5976;
	end
assign N6667 = x_reg_L1_22__retimed_I4004_QOUT;
assign N10416 = !N6667;
assign N10417 = !N10416;
reg x_reg_L1_22__retimed_I4002_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I4002_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22];
	end
assign N6640 = x_reg_L1_22__retimed_I4002_QOUT;
reg x_reg_L1_17__retimed_I3998_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3998_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17];
	end
assign N6631 = x_reg_L1_17__retimed_I3998_QOUT;
reg x_reg_L1_16__retimed_I3994_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3994_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16];
	end
assign N6622 = x_reg_L1_16__retimed_I3994_QOUT;
reg x_reg_L1_14__retimed_I3990_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I3990_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14];
	end
assign N6613 = x_reg_L1_14__retimed_I3990_QOUT;
reg x_reg_L1_13__retimed_I3986_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3986_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13];
	end
assign N6604 = x_reg_L1_13__retimed_I3986_QOUT;
reg x_reg_L1_12__retimed_I3982_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3982_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12];
	end
assign N6595 = x_reg_L1_12__retimed_I3982_QOUT;
reg x_reg_L1_11__retimed_I3978_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I3978_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11];
	end
assign N6586 = x_reg_L1_11__retimed_I3978_QOUT;
reg x_reg_L1_10__retimed_I3974_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I3974_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10];
	end
assign N6577 = x_reg_L1_10__retimed_I3974_QOUT;
reg x_reg_L1_9__retimed_I3970_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I3970_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9];
	end
assign N6568 = x_reg_L1_9__retimed_I3970_QOUT;
reg x_reg_L1_8__retimed_I3966_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3966_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8];
	end
assign N6559 = x_reg_L1_8__retimed_I3966_QOUT;
reg x_reg_L1_7__retimed_I3962_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3962_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7];
	end
assign N6550 = x_reg_L1_7__retimed_I3962_QOUT;
reg x_reg_L1_6__retimed_I3958_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3958_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6];
	end
assign N6541 = x_reg_L1_6__retimed_I3958_QOUT;
reg x_reg_L1_5__retimed_I3954_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3954_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5];
	end
assign N6532 = x_reg_L1_5__retimed_I3954_QOUT;
reg x_reg_L1_4__retimed_I3950_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3950_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4];
	end
assign N6523 = x_reg_L1_4__retimed_I3950_QOUT;
reg x_reg_L1_3__retimed_I3946_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3946_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3];
	end
assign N6514 = x_reg_L1_3__retimed_I3946_QOUT;
reg x_reg_L1_2__retimed_I3942_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3942_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2];
	end
assign N6505 = x_reg_L1_2__retimed_I3942_QOUT;
reg x_reg_L1_1__retimed_I3938_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3938_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1];
	end
assign N6496 = x_reg_L1_1__retimed_I3938_QOUT;
reg x_reg_L1_0__retimed_I3934_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3934_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0];
	end
assign N6487 = x_reg_L1_0__retimed_I3934_QOUT;
reg x_reg_L1_21__retimed_I3930_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I3930_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21];
	end
assign N6478 = x_reg_L1_21__retimed_I3930_QOUT;
reg x_reg_L1_20__retimed_I3926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I3926_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20];
	end
assign N6469 = x_reg_L1_20__retimed_I3926_QOUT;
reg x_reg_L1_19__retimed_I3922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3922_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19];
	end
assign N6460 = x_reg_L1_19__retimed_I3922_QOUT;
reg x_reg_L1_18__retimed_I3918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3918_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18];
	end
assign N6451 = x_reg_L1_18__retimed_I3918_QOUT;
reg x_reg_L1_15__retimed_I3914_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3914_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15];
	end
assign N6442 = x_reg_L1_15__retimed_I3914_QOUT;
reg x_reg_L1_15__retimed_I3911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3911_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70;
	end
assign N6436 = x_reg_L1_15__retimed_I3911_QOUT;
assign N10418 = !N6436;
assign N10419 = !N10418;
reg x_reg_L0_23__retimed_I3863_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3863_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650;
	end
assign N6316 = x_reg_L0_23__retimed_I3863_QOUT;
reg x_reg_L0_22__retimed_I3861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3861_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111;
	end
assign N6311 = x_reg_L0_22__retimed_I3861_QOUT;
reg x_reg_L1_18__retimed_I3854_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3854_QOUT <= N5548;
	end
assign N6227 = x_reg_L1_18__retimed_I3854_QOUT;
reg x_reg_L1_19__retimed_I3851_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3851_QOUT <= N5541;
	end
assign N6220 = x_reg_L1_19__retimed_I3851_QOUT;
reg x_reg_L1_20__retimed_I3848_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I3848_QOUT <= N5534;
	end
assign N6213 = x_reg_L1_20__retimed_I3848_QOUT;
reg x_reg_L1_21__retimed_I3845_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I3845_QOUT <= N5527;
	end
assign N6206 = x_reg_L1_21__retimed_I3845_QOUT;
reg x_reg_L1_23__retimed_I3842_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3842_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0];
	end
assign N6199 = x_reg_L1_23__retimed_I3842_QOUT;
reg x_reg_L1_23__retimed_I3841_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3841_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785;
	end
assign N6197 = x_reg_L1_23__retimed_I3841_QOUT;
reg x_reg_L1_24__retimed_I3838_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I3838_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1];
	end
assign N6190 = x_reg_L1_24__retimed_I3838_QOUT;
reg x_reg_L1_25__retimed_I3835_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I3835_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2];
	end
assign N6183 = x_reg_L1_25__retimed_I3835_QOUT;
reg x_reg_L1_26__retimed_I3832_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I3832_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3];
	end
assign N6176 = x_reg_L1_26__retimed_I3832_QOUT;
reg x_reg_L1_29__retimed_I3824_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I3824_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068;
	end
assign N6157 = x_reg_L1_29__retimed_I3824_QOUT;
reg x_reg_L1_15__retimed_I3818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3818_QOUT <= N5679;
	end
assign N6143 = x_reg_L1_15__retimed_I3818_QOUT;
reg x_reg_L1_0__retimed_I3815_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3815_QOUT <= N5667;
	end
assign N6136 = x_reg_L1_0__retimed_I3815_QOUT;
reg x_reg_L1_1__retimed_I3812_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3812_QOUT <= N5660;
	end
assign N6129 = x_reg_L1_1__retimed_I3812_QOUT;
reg x_reg_L1_2__retimed_I3809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3809_QOUT <= N5653;
	end
assign N6122 = x_reg_L1_2__retimed_I3809_QOUT;
reg x_reg_L1_3__retimed_I3806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3806_QOUT <= N5646;
	end
assign N6115 = x_reg_L1_3__retimed_I3806_QOUT;
reg x_reg_L1_4__retimed_I3803_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3803_QOUT <= N5639;
	end
assign N6108 = x_reg_L1_4__retimed_I3803_QOUT;
reg x_reg_L1_5__retimed_I3800_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3800_QOUT <= N5632;
	end
assign N6101 = x_reg_L1_5__retimed_I3800_QOUT;
reg x_reg_L1_6__retimed_I3797_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3797_QOUT <= N5625;
	end
assign N6094 = x_reg_L1_6__retimed_I3797_QOUT;
reg x_reg_L1_7__retimed_I3794_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3794_QOUT <= N5618;
	end
assign N6087 = x_reg_L1_7__retimed_I3794_QOUT;
reg x_reg_L1_8__retimed_I3791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3791_QOUT <= N5611;
	end
assign N6080 = x_reg_L1_8__retimed_I3791_QOUT;
reg x_reg_L1_9__retimed_I3788_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I3788_QOUT <= N5604;
	end
assign N6073 = x_reg_L1_9__retimed_I3788_QOUT;
reg x_reg_L1_10__retimed_I3785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I3785_QOUT <= N5597;
	end
assign N6066 = x_reg_L1_10__retimed_I3785_QOUT;
reg x_reg_L1_11__retimed_I3782_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I3782_QOUT <= N5590;
	end
assign N6059 = x_reg_L1_11__retimed_I3782_QOUT;
reg x_reg_L1_12__retimed_I3779_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3779_QOUT <= N5583;
	end
assign N6052 = x_reg_L1_12__retimed_I3779_QOUT;
reg x_reg_L1_13__retimed_I3776_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3776_QOUT <= N5576;
	end
assign N6045 = x_reg_L1_13__retimed_I3776_QOUT;
reg x_reg_L1_14__retimed_I3773_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I3773_QOUT <= N5569;
	end
assign N6038 = x_reg_L1_14__retimed_I3773_QOUT;
reg x_reg_L1_16__retimed_I3770_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3770_QOUT <= N5562;
	end
assign N6031 = x_reg_L1_16__retimed_I3770_QOUT;
reg x_reg_L1_17__retimed_I3767_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3767_QOUT <= N5555;
	end
assign N6024 = x_reg_L1_17__retimed_I3767_QOUT;
reg x_reg_L0_31__retimed_I3764_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3764_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6;
	end
assign N6017 = x_reg_L0_31__retimed_I3764_QOUT;
reg x_reg_L0_31__retimed_I3763_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3763_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
	end
assign N6015 = x_reg_L0_31__retimed_I3763_QOUT;
reg x_reg_L0_23__retimed_I3755_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3755_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17;
	end
assign N5991 = x_reg_L0_23__retimed_I3755_QOUT;
reg x_reg_L0_23__retimed_I3754_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3754_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12;
	end
assign N5989 = x_reg_L0_23__retimed_I3754_QOUT;
reg x_reg_L0_15__retimed_I3752_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I3752_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
	end
assign N5976 = x_reg_L0_15__retimed_I3752_QOUT;
reg x_reg_L0_31__retimed_I3657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3657_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282;
	end
assign N5740 = x_reg_L0_31__retimed_I3657_QOUT;
reg x_reg_L0_31__retimed_I3656_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3656_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291;
	end
assign N5738 = x_reg_L0_31__retimed_I3656_QOUT;
reg x_reg_L0_15__retimed_I3631_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I3631_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15];
	end
assign N5679 = x_reg_L0_15__retimed_I3631_QOUT;
reg x_reg_L0_0__retimed_I3626_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I3626_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0];
	end
assign N5667 = x_reg_L0_0__retimed_I3626_QOUT;
reg x_reg_L0_1__retimed_I3623_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I3623_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1];
	end
assign N5660 = x_reg_L0_1__retimed_I3623_QOUT;
reg x_reg_L0_2__retimed_I3620_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I3620_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2];
	end
assign N5653 = x_reg_L0_2__retimed_I3620_QOUT;
reg x_reg_L0_3__retimed_I3617_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I3617_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3];
	end
assign N5646 = x_reg_L0_3__retimed_I3617_QOUT;
reg x_reg_L0_4__retimed_I3614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I3614_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4];
	end
assign N5639 = x_reg_L0_4__retimed_I3614_QOUT;
reg x_reg_L0_5__retimed_I3611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I3611_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5];
	end
assign N5632 = x_reg_L0_5__retimed_I3611_QOUT;
reg x_reg_L0_6__retimed_I3608_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I3608_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6];
	end
assign N5625 = x_reg_L0_6__retimed_I3608_QOUT;
reg x_reg_L0_7__retimed_I3605_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I3605_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7];
	end
assign N5618 = x_reg_L0_7__retimed_I3605_QOUT;
reg x_reg_L0_8__retimed_I3602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I3602_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8];
	end
assign N5611 = x_reg_L0_8__retimed_I3602_QOUT;
reg x_reg_L0_9__retimed_I3599_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I3599_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9];
	end
assign N5604 = x_reg_L0_9__retimed_I3599_QOUT;
reg x_reg_L0_10__retimed_I3596_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I3596_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10];
	end
assign N5597 = x_reg_L0_10__retimed_I3596_QOUT;
reg x_reg_L0_11__retimed_I3593_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I3593_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11];
	end
assign N5590 = x_reg_L0_11__retimed_I3593_QOUT;
reg x_reg_L0_12__retimed_I3590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I3590_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12];
	end
assign N5583 = x_reg_L0_12__retimed_I3590_QOUT;
reg x_reg_L0_13__retimed_I3587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I3587_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13];
	end
assign N5576 = x_reg_L0_13__retimed_I3587_QOUT;
reg x_reg_L0_14__retimed_I3584_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I3584_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14];
	end
assign N5569 = x_reg_L0_14__retimed_I3584_QOUT;
reg x_reg_L0_16__retimed_I3581_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I3581_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16];
	end
assign N5562 = x_reg_L0_16__retimed_I3581_QOUT;
reg x_reg_L0_17__retimed_I3578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I3578_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17];
	end
assign N5555 = x_reg_L0_17__retimed_I3578_QOUT;
reg x_reg_L0_18__retimed_I3575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I3575_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18];
	end
assign N5548 = x_reg_L0_18__retimed_I3575_QOUT;
reg x_reg_L0_19__retimed_I3572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I3572_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19];
	end
assign N5541 = x_reg_L0_19__retimed_I3572_QOUT;
reg x_reg_L0_20__retimed_I3569_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I3569_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20];
	end
assign N5534 = x_reg_L0_20__retimed_I3569_QOUT;
reg x_reg_L0_21__retimed_I3566_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I3566_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21];
	end
assign N5527 = x_reg_L0_21__retimed_I3566_QOUT;
assign bdw_enable = !astall;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132 = !(a_exp[0] & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834 = !((a_exp[7] & a_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172 = !(((a_man[0] | a_man[1]) | a_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155 = !(a_man[10] | a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174 = !(a_man[6] | a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163 = !(a_man[8] | a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183 = !(a_man[4] | a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221 = !(((b_exp[5] & b_exp[4]) & b_exp[7]) & b_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559 = !b_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218 = !(((b_exp[0] & b_exp[1]) & b_exp[2]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249 = !(((b_man[0] | b_man[1]) | b_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232 = !(b_man[10] | b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251 = !(b_man[6] | b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240 = !(b_man[8] | b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260 = !(b_man[4] | b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25] = a_sign ^ b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563 = !b_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408 = a_exp[7] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562 = !b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376 = a_exp[6] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561 = !b_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418 = a_exp[5] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560 = !b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386 = a_exp[4] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360 = a_exp[3] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558 = !b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396 = a_exp[2] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733 = !a_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557 = !b_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557) & a_exp[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 = !b_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404 = !(a_exp[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372 = a_exp[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380 = !(a_exp[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377 = a_exp[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417 = a_exp[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382 = a_exp[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357 = a_exp[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393 = !(a_exp[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 | a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520 = !a_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538 = b_man[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607 = !a_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489 = !(b_man[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541 = !a_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542 = !(b_man[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473 = !a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593 = !(b_man[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561 = !a_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496 = !(b_man[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494 = !a_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548 = !(b_man[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578 = !a_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600 = !(b_man[16] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552 = !a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559 = !(b_man[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484 = !a_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613 = !(b_man[10] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570 = !a_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514 = !(b_man[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516 = !a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502 = !(b_man[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598 = !a_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555 = !(b_man[14] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531 = !a_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605 = !(b_man[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468 = !a_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509 = !(b_man[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507 = !a_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566 = !(b_man[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588 = !a_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467 = !(b_man[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524 = !a_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518 = !(b_man[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610 = !a_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569 = !(b_man[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543 = !a_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471 = !(b_man[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478 = !a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523 = !(b_man[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564 = !a_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575 = !(b_man[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504 = !b_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497 = !a_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477 = !(b_man[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512 = !(b_man[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590 = !(((a_man[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609 = !(b_man[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557 = !(b_man[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506 = !(b_man[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603 = !(b_man[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551 = !(b_man[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500 = !(b_man[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597 = !(b_man[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546 = !(b_man[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493 = !(b_man[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591 = !(b_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540 = !(b_man[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487 = !(b_man[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587 = !(b_man[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534 = !(b_man[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482 = !(b_man[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581 = !(b_man[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528 = !(b_man[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476 = !(b_man[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574 = !(b_man[20] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522 = !(b_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538) | (b_man[22] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340 = ((b_exp[7] | b_exp[5]) | b_exp[6]) | b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336 = ((b_exp[0] | b_exp[1]) | b_exp[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0] = a_exp[0] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565 = a_exp[0] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763 = !((N9273 & N9469) | N9467);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763) & (!N9459)) | (!N9457);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687 & N9195) | N9320);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684 ^ N9187;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687) ^ N9195;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827 = !N10015;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674 = !N9982;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714 & N9390) | N9388);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701) & (!N9329)) | (!N9327);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708) ^ N9122;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701 ^ N9203;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840) & (!N9336)) | (!N9334);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646) ^ N9166;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840 ^ N9219;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763) & (!N9418)) | (!N9416);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838 & N9227) | N9341);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781 ^ N9211;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838) ^ N9227;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737 & N9439) | N9437);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822 = !(((N9374 | N9372) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691) & N9370);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775 = !(N9144 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775 ^ N8595;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822) ^ N9144;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691) & (!N9374)) | (!N9380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650 & N9151) | N9294);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803 ^ N9114;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650) ^ N9151;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724 & N9180) | N9313);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830 ^ N9158;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724) ^ N9180;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750) & (!N9398)) | (!N9396);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677 & N9173) | N9301);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657 ^ N9129;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677) ^ N9173;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773 = !N9985;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820 = !N9988;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667 = !((N9273 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667) & (!N9357)) | (!N9355);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835) ^ N9235;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667 ^ N9259;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] = (!N9281) ^ N9283;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2] = N9289 ^ N9291;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770 = !((N9273 & N9275) | N9362);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770 ^ N9267;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4] = (!N9273) ^ N9275;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793 & N9251) | N9348);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808 ^ N9243;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793) ^ N9251;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919 = (!N7148) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] = (!N10010) ^ N10012;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | (!N8377));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | N8377);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N8377);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439 & N8377;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43 = (N8595 & N8599) | ((!N8595) & N8597);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 & a_sign) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32) & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655 = !(N8357 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & N8357) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633 = N8072 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636 = !(((N7908 | N7910) | N7912) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639 = !(N7934 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53)) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951 = N7159 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941 = !(N7159 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909 = !(N7148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[2]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2]};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946 = N7114 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[3]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913 = (!N7096) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946) | (!(N7114 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917)) | ((!N7096) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[4]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938 = N7088 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938) | (!(N7088 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932) ^ N6921;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905 = ((!N6921) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932)) | ((!N7076) & (!N7078));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6] = (!N9489) ^ N7029;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722 = ((N6183 | N9493) | N9501) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905 & N6915) | (!(N7058 | N7060)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7] = (!N9497) ^ N7050;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950 = ((!N9497) & (!N7050)) | ((!N7066) & (!N7044));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8] = (!N7044) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997 & N6959);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62 = !(N6946 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9] = N7044 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020 = !(((N6962 | N6964) | N6966) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074 | (!N6667));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092 = !(rm[0] & rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 = !(rm[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70 = N6311 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 = !(N10417 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & N6640));
assign x[22] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[21]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & N6478));
assign x[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6206);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[20]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & N6469));
assign x[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6213);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[19]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & N6460));
assign x[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6220);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[18]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & N6451));
assign x[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6227);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[17]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6631));
assign x[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6024);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[16]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6622));
assign x[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6031);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[15]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6442));
assign x[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6143);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[14]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6613));
assign x[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6038);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[13]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6604));
assign x[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6045);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[12]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6595));
assign x[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6052);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[11]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6586));
assign x[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6059);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[10]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6577));
assign x[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6066);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[9]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6568));
assign x[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6073);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[8]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6559));
assign x[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6080);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[7]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6550));
assign x[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6087);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[6]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6541));
assign x[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6094);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[5]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6532));
assign x[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6101);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[4]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6523));
assign x[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6108);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[3]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6514));
assign x[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6115);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6505));
assign x[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6122);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6496));
assign x[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6129);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[0]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & N10419) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & N6487));
assign x[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N6136);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068 = ((N5989 | N5991) | N5976) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074;
assign x[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6157) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]);
assign x[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6157) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]);
assign x[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6157) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & N9501);
assign x[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6157) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & N9493);
assign x[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6157) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & N6176);
assign x[25] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6157) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & N6183);
assign x[24] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6157) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & N6190);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651 = N6316 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0] = ((N5989 | N5991) | N5976) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651;
assign x[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & N6199) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & N6197);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895 = a_sign | b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6) | (a_sign & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_sign) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] & N6017) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]) & N6015);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[31] = (N5738 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285) | ((!N5738) & N5740);
reg x_reg_L1_31__I1187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I1187_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[31];
	end
assign x[31] = x_reg_L1_31__I1187_QOUT;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[0] = x[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[1] = x[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[2] = x[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[3] = x[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[4] = x[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[5] = x[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[6] = x[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[7] = x[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[8] = x[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[9] = x[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[10] = x[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[11] = x[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[12] = x[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[13] = x[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[14] = x[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[15] = x[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[16] = x[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[17] = x[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[18] = x[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[19] = x[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[20] = x[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[21] = x[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[22] = x[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[23] = x[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[24] = x[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[25] = x[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[26] = x[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[27] = x[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[28] = x[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[29] = x[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[30] = x[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[28] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  uLj1TA/ZrR4= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



