/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:10:52 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_1_0 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__30,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42;
wire [15:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51;
wire [24:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3127,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3163,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3169,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3173,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3418,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3525,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3542,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3544,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3554,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3575,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3591,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3604,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3628,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3630,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3644,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3659,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3676,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3710,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3762,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3774,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4152,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4153,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4155,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4163,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4164,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4168,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4171,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4173,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4175,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4178,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4180,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4181,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4186,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4187,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4191,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4193,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4196,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4201,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4204,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4205,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4208,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4212,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4213,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4215,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4221,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4224,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4226,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4228,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4229,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4230,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4231,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4232,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4238,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4239,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4242,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4245,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4254,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4255,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4262,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4264,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4269,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4272,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4274,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4275,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4277,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4278,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4281,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4282,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4287,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4291,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4293,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4296,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4298,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4301,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4304,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4305,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4306,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4310,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4311,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4312,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4313,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4316,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4317,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4319,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4321,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4322,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4323,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4329,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4334,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4336,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4337,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4339,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4340,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4346,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4347,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4351,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4352,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4353,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4356,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4358,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4360,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4361,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4362,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4364,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4365,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4366,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4367,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4368,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4369,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4370,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4371,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4373,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4374,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4375,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4376,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4379,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4380,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4381,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4383,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4385,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4386,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4388,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4391,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4393,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4396,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4397,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4398,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4400,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4401,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4403,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4405,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4410,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4418,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4420,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4423,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4425,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4429,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4434,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4440,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4441,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4443,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4445,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4447,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4460,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4461,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4462,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4463,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4465,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4472,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4476,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4495,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4506,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4513,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4515,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4518,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4520,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4521,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4522,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4524,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4525,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4526,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4527,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4528,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4530,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4532,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4536,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4537,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4538,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4539,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4541,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4542,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4543,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4544,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4546,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4547,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4549,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4552,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4554,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4559,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4560,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4564,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4566,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4569,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4571,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4580,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4585,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4586,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4591,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4595,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4597,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4602,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4605,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4607,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4618,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4622,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4623,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4628,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4635,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4639,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4640,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4641,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4646,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4647,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4649,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4654,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4659,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4660,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4663,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4665,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4667,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4669,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4671,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4672,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4673,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4676,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4677,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4678,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4681,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4682,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4685,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4687,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4688,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4689,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4694,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4697,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4700,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4701,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4702,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4707,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4709,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4711,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4712,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4713,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4715,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4716,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4720,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4722,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4723,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4724,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4727,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4728,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4729,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4732,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4733,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4734,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4735,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4738,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4742,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4743,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4744,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4746,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4749,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4750,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4752,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4753,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4755,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4756,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4758,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4761,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4763,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4764,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4765,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4770,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4771,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4773,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4776,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4778,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4779,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4780,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4782,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4791,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4792,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4793,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4796,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4797,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4798,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4799,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4800,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4803,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4804,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4806,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4807,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4808,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4809,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4810,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4812,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4813,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4814,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4815,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4816,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4817,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4819,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4821,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4823,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4824,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4825,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4828,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4829,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4830,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4831,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4833,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4834,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4836,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4839,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4841,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4843,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4844,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4845,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4846,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4847,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4848,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4850,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4851,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4854,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4857,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4858,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4859,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4860,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4861,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4862,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4865,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4867,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4868,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4871,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4872,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4876,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4878,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4881,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4882,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4883,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4884,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4885,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4886,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4887,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4888,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4889,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4890,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4891,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4892,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4895,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4898,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4899,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4901,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4902,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4905,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4906,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4907,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4908,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4909,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4910,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4912,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4913,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4914,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4916,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4919,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4920,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4922,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4923,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4924,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4925,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4926,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4927,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4928,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4930,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4931,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4932,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4933,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4936,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4937,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4938,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4941,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4942,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4944,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4945,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4947,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4949,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4950,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4951,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4952,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4954,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4955,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4956,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4957,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4961,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4962,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4963,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4965,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4966,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4970,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4972,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4974,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4975,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4977,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4978,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4979,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4980,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4982,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4983,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4984,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4985,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4986,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4987,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4989,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4990,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4991,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4993,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4994,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4996,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4997,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5000,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5001,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5002,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5005,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5006,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5007,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5009,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5012,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5013,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5014,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5016,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5017,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5018,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5019,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5021,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5024,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5025,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5026,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5027,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5028,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5029,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5030,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5031,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5032,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5035,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5036,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5037,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5039,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5040,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5041,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5042,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5043,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5047,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5050,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5051,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5052,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5053,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5054,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5055,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5056,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5057,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5058,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5059,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5060,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5063,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5068,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5070,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5082,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5098,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5103,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5107,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5109,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5111,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5117,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5119,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5126,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5128,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5136,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5138,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5160,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6178,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6191,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6200,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6207,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6231,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6238,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6239,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6269,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6274,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6277,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6279,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6311,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6319,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6321,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6323,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6334,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6336,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6351,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6353,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6355,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6379,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6381,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6383,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6385,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6393,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6397,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6409,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6423,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6431,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6438,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6440,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6476,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6505,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6832,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6833,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6834,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6835,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6837,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6839,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6840,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6841,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6842,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6843,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6844,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6845,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6846,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6847,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6848,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6849,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6850,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6851,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6852,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6853,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6854,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6856,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6857,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6859,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6860,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6861,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6863,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6864,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6865,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6866,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6868,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6869,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6870,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6871,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6873,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6874,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6875,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6876,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6877,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6878,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6880,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6881,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6882,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6883,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6884,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6886,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6887,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6888,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6889,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6891,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6892,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6893,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6894,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6895,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6896,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6897,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6899,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6900,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6901,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6902,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6903,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6904,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6905,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6907,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6908,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6909,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6910,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6911,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6912,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6913,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6914,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6916,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6917,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6918,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6919,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6920,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6921,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6922,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6923,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6924,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6925,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6927,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6929,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6931,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6932,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6933,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6935,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6936,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6937,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6939,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6940,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6941,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6943,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6944,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6945,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6946,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6948,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6949,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6950,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6951,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6953,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6954,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6955,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6956,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6957,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6958,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6960,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6961,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6962,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6963,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6964,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6965,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6966,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6968,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6969,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6970,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6971,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6972,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6974,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6975,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6976,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6977,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6978,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6981,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6982,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6985,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6986,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6987,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6988,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6989,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6990,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6992,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6994,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6995,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6996,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6997,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6999,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7000,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7001,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7002,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7003,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7004,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7005,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7006,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7007,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7009,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7010,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7011,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7012,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7013,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7014,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7015,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7018,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7019,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7020,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7021,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7022,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7023,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7025,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7026,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7028,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7029,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7031,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7032,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7034,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7035,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7036,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7037,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7038,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7039,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7040,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7043,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7044,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7045,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7046,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7047,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7048,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7049,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7051,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7052,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7054,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7055,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7056,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7057,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7058,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7060,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7061,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7063,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7064,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7065,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7066,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7068,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7069,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7071,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7072,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7073,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7074,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7075,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7077,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7078,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7079,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7080,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7081,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7082,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7083,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7084,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7086,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7087,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7088,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7089,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7091,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7093,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7094,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7095,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7097,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7098,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7101,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7102,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7103,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7104,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7105,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7106,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7107,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7110,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7111,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7112,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7113,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7114,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7115,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7116,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7117,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7118,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7120,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7121,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7122,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7123,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7127,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7128,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7129,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7130,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7132,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7133,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7135,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7136,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7137,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7138,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7141,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7143,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7145,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7152,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7153,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7154,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7155,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7160,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7162,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7164,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7166,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7169,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7171,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7173,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7174,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7175,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7178,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7180,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7181,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7184,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7187,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7188,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7191,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7193,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7194,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7196,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7197,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7200,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7204,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7205,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7208,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7212,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7215,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7219,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7221,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7224,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7228,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7229,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7232,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7236,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7238,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7245,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7248,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7249,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7253,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7254,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7255,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7261,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7264,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7269,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7270,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7271,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7272,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7274,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7275,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7276,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7277,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7279,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7281,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7282,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7283,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7287,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7289,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7290,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7291,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7293,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7294,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7296,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7298,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7300,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7301,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7302,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7303,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7305,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7306,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7308,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7309,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7311,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7312,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7313,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7316,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7317,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7319,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7322,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7323,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7325,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7331,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7334,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7336,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7337,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7340,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7342,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7345,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7346,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7347,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7351,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7352,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7353,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7356,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7357,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7358,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7359,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7360,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7362,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7365,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7366,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7367,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7368,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7369,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7370,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7371,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7372,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7373,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7374,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7375,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7376,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7378,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7379,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7380,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7381,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7382,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7383,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7384,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7385,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7386,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7387,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7388,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7389,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7390,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7391,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7396,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7398,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7401,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7405,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7406,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7408,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7409,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7410,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7418,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7423,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7429,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7431,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7432,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7435,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7440,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7441,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7445,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7459,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7460,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7463,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7469,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7472,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7475,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7495,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7502,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7505,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7506,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7513,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7516,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7517,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7518,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7519,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7520,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7522,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7524,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7526,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7527,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7529,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7530,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7531,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7534,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7535,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7536,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7538,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7539,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7541,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7542,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7544,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7545,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7547,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7551,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7554,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7555,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7559,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7560,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7561,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7566,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7567,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7573,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7575,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7577,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7578,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7580,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7582,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7587,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7589,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7591,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7595,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7602,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7604,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7607,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7609,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7611,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7613,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7614,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7622,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7625,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7630,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7633,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7639,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7640,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7641,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7644,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7646,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7647,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7650,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7652,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7655,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7656,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7658,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7659,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7660,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7665,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7666,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7669,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7672,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7673,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7676,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7677,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7679,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7681,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7682,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7684,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7685,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7689,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7693,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7694,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7697,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7699,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7700,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7702,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7706,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7707,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7710,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7711,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7712,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8572,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8575,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8586,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8589,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8602,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8604,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8605,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8607,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8625,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8639,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8651,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8655,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8665,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8671,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8677,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8707,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8715,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8718,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8720,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8731,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8733,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8734,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8736,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8743,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8745,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8746,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8747,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8750,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8752,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8756,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8762,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8768,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8769,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8770,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8774,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8777,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8792,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8793,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8795,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8796,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8803,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8806,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8814,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8817,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8822,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8830,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8831,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8835,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8836,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8839,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8840,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8843,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8846,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8848,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8854,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8861,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8862,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8863,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8866,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8867,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8868,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8873,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8879,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8881,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8892,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8893,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8898,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8901,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8909,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8911,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8913,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8925,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8926,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8928,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8929,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8930,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8931,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8940,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8942,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8944,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8946,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8949,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8953,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8956,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8967,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8970,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8971,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8980,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8983,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8989,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8994,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8999,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9003,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9004,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9006,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9008,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9010,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9014,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9015,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9026,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9029,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9030,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9034,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9035,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9038,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9039,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9040,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9042,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9054,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9056,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9059,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9065,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9068,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9070,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9080,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9081,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9086,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9087,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9088,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9098,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9110,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9112,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9126,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9128,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9129,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9130,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9172,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9174,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9195,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9207,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9218,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9221,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9231,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9236,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9242,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9248,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9282,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9283,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9294,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13732,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13738,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13813,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13851,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26089,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26095,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26111,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26143,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26168,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26200,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26213,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26219,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26229,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26230,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26236,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26253,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26312,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26314,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26322,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26325,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26340,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26352,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26359,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26461,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26561,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26585,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26587,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26611,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26688,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26710,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26737;
wire N12256,N12258,N12260,N12465,N12467,N12472,N12474 
	,N12479,N12481,N12486,N12488,N12493,N12495,N12500,N12502 
	,N12528,N12530,N12535,N12537,N12544,N12547,N12549,N12554 
	,N12569,N12574,N12682,N12687,N12712,N12719,N12722,N12729 
	,N12734,N12737,N12739,N12742,N12744,N12747,N12749,N12752 
	,N12754,N12834,N12863,N12894,N12896,N12942,N12967,N12969 
	,N12983,N12990,N13013,N13023,N13035,N13068,N13070,N13072 
	,N13106,N13108,N13125,N13132,N13134,N13138,N13142,N13146 
	,N13456,N13460,N13643,N13644,N13645,N13646,N13647,N13648 
	,N13649,N13650;
reg x_reg_8__retimed_I7925_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I7925_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9284;
	end
assign N13460 = x_reg_8__retimed_I7925_QOUT;
reg x_reg_10__retimed_I7923_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I7923_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9247;
	end
assign N13456 = x_reg_10__retimed_I7923_QOUT;
reg x_reg_2__retimed_I7820_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7820_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9038;
	end
assign N13146 = x_reg_2__retimed_I7820_QOUT;
reg x_reg_18__retimed_I7818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7818_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8949;
	end
assign N13142 = x_reg_18__retimed_I7818_QOUT;
reg x_reg_15__retimed_I7816_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7816_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8839;
	end
assign N13138 = x_reg_15__retimed_I7816_QOUT;
reg x_reg_15__retimed_I7814_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7814_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8750;
	end
assign N13134 = x_reg_15__retimed_I7814_QOUT;
reg x_reg_2__retimed_I7813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7813_QOUT <= N13125;
	end
assign N13132 = x_reg_2__retimed_I7813_QOUT;
reg x_reg_15__retimed_I7802_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7802_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209;
	end
assign N13108 = x_reg_15__retimed_I7802_QOUT;
reg x_reg_15__retimed_I7801_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7801_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805;
	end
assign N13106 = x_reg_15__retimed_I7801_QOUT;
reg x_reg_2__retimed_I7790_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7790_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26553;
	end
assign N13072 = x_reg_2__retimed_I7790_QOUT;
reg x_reg_2__retimed_I7789_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7789_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26548;
	end
assign N13070 = x_reg_2__retimed_I7789_QOUT;
reg x_reg_2__retimed_I7788_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7788_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8944;
	end
assign N13068 = x_reg_2__retimed_I7788_QOUT;
reg x_reg_15__retimed_I7775_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7775_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922;
	end
assign N13035 = x_reg_15__retimed_I7775_QOUT;
reg x_reg_2__retimed_I7771_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7771_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206;
	end
assign N13023 = x_reg_2__retimed_I7771_QOUT;
reg x_reg_2__retimed_I7767_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7767_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26565;
	end
assign N13013 = x_reg_2__retimed_I7767_QOUT;
reg x_reg_11__retimed_I7760_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I7760_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103;
	end
assign N12990 = x_reg_11__retimed_I7760_QOUT;
reg x_reg_18__retimed_I7758_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7758_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013;
	end
assign N12983 = x_reg_18__retimed_I7758_QOUT;
reg x_reg_11__retimed_I7754_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I7754_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8983;
	end
assign N12969 = x_reg_11__retimed_I7754_QOUT;
reg x_reg_11__retimed_I7753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I7753_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8806;
	end
assign N12967 = x_reg_11__retimed_I7753_QOUT;
reg x_reg_10__retimed_I7745_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I7745_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986;
	end
assign N12942 = x_reg_10__retimed_I7745_QOUT;
reg x_reg_15__retimed_I7730_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7730_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156;
	end
assign N12896 = x_reg_15__retimed_I7730_QOUT;
reg x_reg_15__retimed_I7729_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7729_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993;
	end
assign N12894 = x_reg_15__retimed_I7729_QOUT;
reg x_reg_9__retimed_I7718_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I7718_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071;
	end
assign N12863 = x_reg_9__retimed_I7718_QOUT;
reg x_reg_10__retimed_I7708_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I7708_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9065;
	end
assign N12834 = x_reg_10__retimed_I7708_QOUT;
reg x_reg_19__retimed_I7678_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I7678_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9030;
	end
assign N12754 = x_reg_19__retimed_I7678_QOUT;
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I8016 (.Y(N13643), .A(N12754));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I8017 (.Y(N13644), .A(N13643));
reg x_reg_19__retimed_I7677_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I7677_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8861;
	end
assign N12752 = x_reg_19__retimed_I7677_QOUT;
reg x_reg_14__retimed_I7676_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I7676_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9174;
	end
assign N12749 = x_reg_14__retimed_I7676_QOUT;
reg x_reg_14__retimed_I7675_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I7675_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8746;
	end
assign N12747 = x_reg_14__retimed_I7675_QOUT;
reg x_reg_1__retimed_I7674_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I7674_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610;
	end
assign N12744 = x_reg_1__retimed_I7674_QOUT;
reg x_reg_1__retimed_I7673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I7673_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772;
	end
assign N12742 = x_reg_1__retimed_I7673_QOUT;
reg x_reg_3__retimed_I7672_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I7672_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262;
	end
assign N12739 = x_reg_3__retimed_I7672_QOUT;
reg x_reg_3__retimed_I7671_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I7671_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686;
	end
assign N12737 = x_reg_3__retimed_I7671_QOUT;
reg x_reg_8__retimed_I7670_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I7670_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075;
	end
assign N12734 = x_reg_8__retimed_I7670_QOUT;
reg x_reg_8__retimed_I7668_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I7668_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239;
	end
assign N12729 = x_reg_8__retimed_I7668_QOUT;
reg x_reg_5__retimed_I7665_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I7665_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578;
	end
assign N12722 = x_reg_5__retimed_I7665_QOUT;
reg x_reg_9__retimed_I7664_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I7664_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917;
	end
assign N12719 = x_reg_9__retimed_I7664_QOUT;
reg x_reg_9__retimed_I7661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I7661_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8956;
	end
assign N12712 = x_reg_9__retimed_I7661_QOUT;
reg x_reg_0__retimed_I7651_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I7651_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8873;
	end
assign N12687 = x_reg_0__retimed_I7651_QOUT;
reg x_reg_0__retimed_I7649_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I7649_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8715;
	end
assign N12682 = x_reg_0__retimed_I7649_QOUT;
reg x_reg_11__retimed_I7609_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I7609_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9259;
	end
assign N12574 = x_reg_11__retimed_I7609_QOUT;
reg x_reg_19__retimed_I7607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I7607_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26692;
	end
assign N12569 = x_reg_19__retimed_I7607_QOUT;
reg x_reg_7__retimed_I7601_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I7601_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8796;
	end
assign N12554 = x_reg_7__retimed_I7601_QOUT;
reg x_reg_15__retimed_I7599_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7599_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170;
	end
assign N12549 = x_reg_15__retimed_I7599_QOUT;
reg x_reg_15__retimed_I7598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7598_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26737;
	end
assign N12547 = x_reg_15__retimed_I7598_QOUT;
reg x_reg_14__retimed_I7597_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I7597_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8879;
	end
assign N12544 = x_reg_14__retimed_I7597_QOUT;
reg x_reg_13__retimed_I7594_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I7594_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9140;
	end
assign N12537 = x_reg_13__retimed_I7594_QOUT;
reg x_reg_13__retimed_I7593_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I7593_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9292;
	end
assign N12535 = x_reg_13__retimed_I7593_QOUT;
reg x_reg_12__retimed_I7591_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I7591_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8651;
	end
assign N12530 = x_reg_12__retimed_I7591_QOUT;
reg x_reg_12__retimed_I7590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I7590_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8803;
	end
assign N12528 = x_reg_12__retimed_I7590_QOUT;
reg x_reg_22__retimed_I7579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7579_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8817;
	end
assign N12502 = x_reg_22__retimed_I7579_QOUT;
reg x_reg_22__retimed_I7578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7578_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8989;
	end
assign N12500 = x_reg_22__retimed_I7578_QOUT;
reg x_reg_21__retimed_I7576_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I7576_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9080;
	end
assign N12495 = x_reg_21__retimed_I7576_QOUT;
reg x_reg_21__retimed_I7575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I7575_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9242;
	end
assign N12493 = x_reg_21__retimed_I7575_QOUT;
reg x_reg_20__retimed_I7573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I7573_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8584;
	end
assign N12488 = x_reg_20__retimed_I7573_QOUT;
reg x_reg_20__retimed_I7572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I7572_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8752;
	end
assign N12486 = x_reg_20__retimed_I7572_QOUT;
reg x_reg_18__retimed_I7570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7570_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8846;
	end
assign N12481 = x_reg_18__retimed_I7570_QOUT;
reg x_reg_18__retimed_I7569_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7569_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9015;
	end
assign N12479 = x_reg_18__retimed_I7569_QOUT;
reg x_reg_17__retimed_I7567_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I7567_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9108;
	end
assign N12474 = x_reg_17__retimed_I7567_QOUT;
reg x_reg_17__retimed_I7566_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I7566_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9265;
	end
assign N12472 = x_reg_17__retimed_I7566_QOUT;
reg x_reg_16__retimed_I7564_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I7564_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8616;
	end
assign N12467 = x_reg_16__retimed_I7564_QOUT;
reg x_reg_16__retimed_I7563_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I7563_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8774;
	end
assign N12465 = x_reg_16__retimed_I7563_QOUT;
reg x_reg_18__retimed_I7472_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7472_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67;
	end
assign N12260 = x_reg_18__retimed_I7472_QOUT;
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I8018 (.Y(N13645), .A(N12260));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I8019 (.Y(N13646), .A(N13645));
reg x_reg_18__retimed_I7471_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7471_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9934;
	end
assign N12258 = x_reg_18__retimed_I7471_QOUT;
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I8020 (.Y(N13647), .A(N12258));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I8021 (.Y(N13648), .A(N13647));
reg x_reg_18__retimed_I7470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7470_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320;
	end
assign N12256 = x_reg_18__retimed_I7470_QOUT;
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I8022 (.Y(N13649), .A(N12256));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I8023 (.Y(N13650), .A(N13649));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I0 (.Y(bdw_enable), .A(astall));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3127), .A(a_exp[6]), .B(a_exp[5]));
AND4XL float_div_cynw_cm_float_rcp_E8_M23_1_I2 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3125), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL float_div_cynw_cm_float_rcp_E8_M23_1_I3 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13813), .A(a_exp[7]), .B(a_exp[0]), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3125));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I4 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3127), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13813));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I5 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I6 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .A(a_man[2]));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_1_I7 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3163), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I8 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3167), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(a_man[0]), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3163), .D(a_man[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I9 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3148), .A(a_man[10]), .B(a_man[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I10 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3169), .A(a_man[6]), .B(a_man[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I11 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3158), .A(a_man[8]), .B(a_man[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I12 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3179), .A(a_man[4]), .B(a_man[3]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_1_I13 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3161), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3148), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3169), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3158), .D(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3179));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_1_I14 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3173), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_1_I15 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3183), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I16 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3167), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3161), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3173), .D(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3183));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I17 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I18 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I19 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3335), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I20 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3326), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I21 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3338), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I22 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3330), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_1_I23 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3328), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3335), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3326), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3338), .D(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3330));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I24 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3328), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I25 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[1]), .A(a_exp[1]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I26 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[0]), .A(a_exp[0]));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I27 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I28 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[1]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I29 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2]), .A(a_exp[2]));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I30 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I31 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3240), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I32 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[3]), .A(a_exp[3]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I33 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3240), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[3]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I34 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[5]), .A(a_exp[5]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I35 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4]), .A(a_exp[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I36 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3256), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I37 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3256), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I38 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3248), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I39 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3248));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_1_I40 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3292), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[3]), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I41 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I42 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[6]), .A(a_exp[6]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I43 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[6]));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I44 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3241), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254));
MXI2XL float_div_cynw_cm_float_rcp_E8_M23_1_I45 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3241), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I46 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3233), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I47 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7]), .A(a_exp[7]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I48 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3244), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3233), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7]));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I49 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I50 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3295), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[7]));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I51 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[0]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I52 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I53 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[1]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[1]));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I54 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3289), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3295), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[0]), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[4]), .D(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[1]));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I55 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[8]), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[6]), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237), .D(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7]));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_1_I56 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__17), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3292), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3289), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[8]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I57 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__30), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__17));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_1_I58 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N447), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9), .A1N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__30));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I59 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N447));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_1_I60 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26688), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]), .D(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I61 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26688));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I62 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9934), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I63 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A(a_man[22]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I64 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A(a_man[21]));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I65 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A(a_man[19]));
CLKINVX4 float_div_cynw_cm_float_rcp_E8_M23_1_I66 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350), .A(a_man[18]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I67 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I68 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(a_man[17]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I69 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I70 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4601), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261), .B(a_man[20]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I71 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A(a_man[20]));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I72 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350));
CLKINVX12 float_div_cynw_cm_float_rcp_E8_M23_1_I73 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015));
CLKINVX8 float_div_cynw_cm_float_rcp_E8_M23_1_I74 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I75 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789));
CLKINVX8 float_div_cynw_cm_float_rcp_E8_M23_1_I76 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .A(a_man[16]));
CLKINVX8 float_div_cynw_cm_float_rcp_E8_M23_1_I77 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I78 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B(a_man[17]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I79 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I80 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I81 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I82 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4246), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4601), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093), .B1(a_man[21]));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I83 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I84 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I85 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516), .A(a_man[17]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I86 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13759), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516));
CLKINVX12 float_div_cynw_cm_float_rcp_E8_M23_1_I87 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13759));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I88 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I89 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I90 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4385), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I91 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4385), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I92 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4821), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I93 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4246), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4821), .B1(a_man[22]));
NOR2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I94 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I95 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I96 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4867), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I97 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4867), .B(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I98 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4979), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I99 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N501), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4979), .B(a_man[22]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N501));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4646), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141), .A(a_man[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4231), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4374), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4646), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4231), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4824), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5025), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4824), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I109 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5042), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4374), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5025), .B1(a_man[21]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I110 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789));
NOR2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I111 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .A(a_man[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_1_I113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4418), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .A1N(a_man[19]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4232), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4600), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4418), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4232), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5042), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4600), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4419), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5029), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4156), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4419), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5029), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4847), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4603), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4803), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4847), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4603), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4817), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4156), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4803), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5041), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4198), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5041), .B0(a_man[19]), .B1(a_man[20]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5030), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4373), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4198), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5030), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4817), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4373), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576));
AOI22X2 float_div_cynw_cm_float_rcp_E8_M23_1_I143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4421), .A0(a_man[16]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4421));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I145 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4199), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4955), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4199), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4225), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4626), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4225), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I161 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I162 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4376), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4581), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4626), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4376), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4596), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4955), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4581), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4816), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I166 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4319), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I167 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4993), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4816), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4319), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I168 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B1(a_man[19]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I169 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I170 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4848), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4808), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4848), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I172 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4155), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4993), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4808), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I173 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N497), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4596), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4155), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I174 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976), .A(1'B1), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N497));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9129), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9129), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8909), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8989), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8909));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8817), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4994), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875), .B1(a_man[19]));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .A(a_man[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22X2 float_div_cynw_cm_float_rcp_E8_M23_1_I196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4713), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(a_man[17]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4713));
CLKINVX8 float_div_cynw_cm_float_rcp_E8_M23_1_I198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .B(a_man[17]));
AOI22X4 float_div_cynw_cm_float_rcp_E8_M23_1_I200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I201 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4585), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4728), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4994), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4585), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I203 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4400), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I207 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4158), .A0(a_man[17]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4358), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4400), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4158), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4369), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4728), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4358), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I213 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958), .A0(a_man[17]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4594), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I215 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .B1(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I216 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5117), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I217 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4770), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4594), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5117), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4631), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4627), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I221 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4586), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4631), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4627), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4954), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4770), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4586), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4369), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4954), .B1(a_man[22]));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .A(a_man[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4334), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4360), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4508), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4334), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4360), .B1(a_man[20]));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
CLKBUFX6 float_div_cynw_cm_float_rcp_E8_M23_1_I229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995));
AO22XL float_div_cynw_cm_float_rcp_E8_M23_1_I230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4180), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4957), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5157), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4180), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4957), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4152), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4508), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5157), .B1(a_man[21]));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4367), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13558), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762));
BUFX3 float_div_cynw_cm_float_rcp_E8_M23_1_I245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13558));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4890), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4546), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4367), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4890), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935), .A0(a_man[17]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4405), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777), .B1(a_man[19]));
AO22XL float_div_cynw_cm_float_rcp_E8_M23_1_I252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4825), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4825));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4401), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4361), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4405), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4401), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4727), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4546), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4361), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N495), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4152), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4727), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I258 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9026), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N495));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I259 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I260 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4495), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5143), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726), .B(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4580), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4495), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5143), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[16]), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4580));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7205), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[16]));
CLKINVX4 float_div_cynw_cm_float_rcp_E8_M23_1_I268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .A(a_man[14]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I269 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4560), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_1_I271 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[17]), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4560), .A1N(a_man[21]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I272 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[17]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I273 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7179), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I274 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .A(a_man[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I275 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7656), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7463), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7205), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7179), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I276 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7595), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[17]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I277 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[33]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[32]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7656), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7595), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5133), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5160), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4292), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5133), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5160), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4980), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4938), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4980), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4952), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4292), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4938), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4149), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I289 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4669), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I290 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4333), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4149), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4669), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I291 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I293 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4183), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4181), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5161), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4183), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4181), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4507), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4333), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5161), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N494), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4952), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4507), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I299 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8631), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9218), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N494), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[32]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I300 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9026), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[33]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8631));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I302 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I303 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7651), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX8 float_div_cynw_cm_float_rcp_E8_M23_1_I304 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .A(a_man[12]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I305 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4532), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4275), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4532), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4920), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4356), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4275), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4920), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I310 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4926), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4494), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4926), .B(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[15]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4356), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4494), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I314 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7710), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I315 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7380), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7188), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7651), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7710));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5115), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5145), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I318 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4274), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5115), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5145), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I319 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4317), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4924), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5069), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4317), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4924), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I323 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4734), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I324 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4691), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4734), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I325 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5156), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5069), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4691), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I326 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339), .A0(a_man[22]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4274), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5156));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I327 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7322), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I328 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7233), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I329 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .A(a_man[11]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I330 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7609), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7415), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7322), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7233), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7680), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I333 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6882), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7573), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7609), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7680), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I334 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[32]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7463), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7380), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6882));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5148), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4906), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5148), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4941), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I340 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5083), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4906), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4941), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4754), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4862), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4709), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4862), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I345 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4724), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5083), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4709), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I346 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4947), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I347 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4445), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I348 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5132), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4947), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4445), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I349 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4982), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I350 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4942), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4982), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I351 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4291), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5132), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4942), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N493), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4724), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4291), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I353 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8814), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8662), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N493), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[31]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I354 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[32]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9218), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8814));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7293), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7261), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6849), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7707), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX8 float_div_cynw_cm_float_rcp_E8_M23_1_I361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .A(a_man[10]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I362 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7451), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7254), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6849), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7707), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I363 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7112), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6917), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7293), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7261), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7451));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6877), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4705), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5001), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4888), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4705), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5001));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4925), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5068), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4888), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4925), .B1(a_man[21]));
AOI22X2 float_div_cynw_cm_float_rcp_E8_M23_1_I370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I371 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5116), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(a_man[17]), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I372 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I373 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4695), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4844), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5116), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4695));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I377 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I378 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4473), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4936), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4844), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4473), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5068), .A1(a_man[22]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4936));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6935), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I382 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6908), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I384 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6950), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7642), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6877), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6935), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6908));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I385 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7498), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7301), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6950), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7415), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6917));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I386 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[31]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7573), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7112), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7498));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I387 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4285), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I388 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I389 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4681), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4285), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I390 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I391 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I392 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4711), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I393 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4860), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4681), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4711), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4528), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4643), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4492), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4528), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4643), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I398 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4506), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4860), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4492), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4245), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4722), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4245), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4223), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4905), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4722), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4223), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4756), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I404 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5112), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4712), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4756), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5112), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5082), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4905), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4712), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N492), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4506), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5082), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I409 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9014), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8843), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N492), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[30]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I410 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[31]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8662), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9014));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8768), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7319), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7290), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX12 float_div_cynw_cm_float_rcp_E8_M23_1_I416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .A(a_man[9]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I417 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6902), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7591), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7319), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7290), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7347), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4889), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I421 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4477), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I422 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4622), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4889), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4477));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I423 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4298), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I424 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4251), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4298), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4707), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4622), .B0(a_man[21]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4251));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4490), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I428 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I429 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4778), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4667), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4490), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4778), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4997), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I432 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4696), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4997), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I433 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4843), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4667), .B0(a_man[21]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4696));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[12]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4707), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4843), .B1(a_man[22]));
CLKBUFX2 float_div_cynw_cm_float_rcp_E8_M23_1_I435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[12]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7435), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7375), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I438 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7285), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7097), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7435), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7375));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I439 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7336), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7147), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7254), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6902), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7285));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I440 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6905), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6874), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX12 float_div_cynw_cm_float_rcp_E8_M23_1_I442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .A(a_man[8]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I443 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6853), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7544), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6905), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6874), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I444 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I445 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7405), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I446 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7676), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7484), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6853), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7405), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7591));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I447 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6840), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7530), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7676), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7642), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7147));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I448 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[30]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7301), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7336), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6840));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I449 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I450 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4482), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4461), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4482), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4497), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4641), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4461), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4497), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I456 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4315), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I458 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I459 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4416), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I460 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4272), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4315), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4416), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I461 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4288), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4641), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4272), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I462 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I463 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I464 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4504), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5019), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4680), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4504), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5019), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4536), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I469 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4886), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I471 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4498), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4536), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4886), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I472 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4859), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4680), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4498), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I473 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N491), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4288), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4859), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I474 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9207), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9039), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N491), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[29]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I475 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8843), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[30]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9207));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I476 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7402), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4444), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I481 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5051), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4176), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4444), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5051));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I485 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4868), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I486 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4530), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I487 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4823), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4868), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4530), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I488 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4269), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4176), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4823), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I489 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I490 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5059), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I491 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4338), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4220), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5059), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4338));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I494 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I495 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4424), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I496 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4549), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I497 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4257), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4424), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4549), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I498 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4396), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4220), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4257), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I499 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[10]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4269), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4396), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I500 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7547), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[10]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I501 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7432), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I502 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7693), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7502), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7402), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7547), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7432));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I503 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I504 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7492), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I505 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7464), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I506 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I507 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4668), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I508 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I509 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4256), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I510 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4397), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4668), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4256));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5091), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4755), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5047), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5091), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4755), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4491), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4397), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5047), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4267), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I517 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4552), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I518 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4443), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4267), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4552), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4772), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I520 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4478), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4772), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4621), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4443), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4478), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I522 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[11]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4491), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4621), .B1(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I523 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I524 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7523), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I525 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7192), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7000), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7492), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7464), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7523));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I526 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7128), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6932), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7693), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7544), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7192));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I527 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7022), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I528 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6990), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I529 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7373), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I530 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7345), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX12 float_div_cynw_cm_float_rcp_E8_M23_1_I531 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .A(a_man[7]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I532 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7307), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7116), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7373), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7345), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I533 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7624), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7431), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7022), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6990), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7307));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I534 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6933), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I535 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7051), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I536 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6961), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I537 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7236), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7048), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6933), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7051), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6961));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6958), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6929), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I540 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .A(a_man[6]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I541 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7370), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7176), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6958), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6929), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I542 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6988), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I543 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I544 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4221), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4830), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I547 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4975), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4221), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4830));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I548 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4647), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I549 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4316), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4602), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4647), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4316), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5063), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4975), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4602), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I552 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4391), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I553 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5138), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I554 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5017), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4391), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5138), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I555 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4205), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I557 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4337), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I558 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5053), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4205), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4337), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I559 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4175), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5017), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5053), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I560 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[9]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5063), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4175), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I561 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7160), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7019), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I563 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6871), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7563), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6988), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7160), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7019));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I564 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7579), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7383), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7116), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7370), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6871));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I565 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7516), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7318), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7431), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7048), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7579));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I566 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7560), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7368), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7484), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7128), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7516));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I567 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7174), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6981), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7624), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7236), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7097));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I568 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[29]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7560), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7174), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7530));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4238), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I571 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I573 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4277), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4415), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4238), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4277), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I575 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I576 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4182), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I577 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5111), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4182), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I578 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I579 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I580 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4196), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I581 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5066), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5111), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4196), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I582 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5080), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4415), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5066), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I583 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510), .A0(a_man[17]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I584 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4284), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I585 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4202), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I587 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4798), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4202), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I588 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4460), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4284), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4798), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I589 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4687), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4321), .A0(a_man[17]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4687), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I592 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4664), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I593 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4278), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4321), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4664), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I594 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4640), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4460), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4278), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N490), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5080), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4640), .B1(a_man[22]));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I596 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[10]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7136), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I598 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7049), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7078), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I600 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7258), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7068), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7136), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7049), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7078));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I601 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7429), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I602 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7399), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX4 float_div_cynw_cm_float_rcp_E8_M23_1_I603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .A(a_man[5]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I604 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7054), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6856), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7429), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7399), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I605 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7107), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I606 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7646), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7454), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7054), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7107), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I607 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7082), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6887), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7502), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7258), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7646));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I608 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7013), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7706), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7082), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6932), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7318));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I609 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[28]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7013), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6981), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7368));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I610 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8648), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9231), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N490), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[28]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I611 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9039), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[29]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8648));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I612 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I613 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8589), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I614 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4636), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I615 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5036), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4636), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I616 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I617 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I618 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5070), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I619 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4193), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5036), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5070), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4885), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4991), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4841), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4885), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4991), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4858), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4193), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4841), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I626 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5077), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I627 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5100), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I629 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4571), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5100), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I630 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4237), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5077), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4571), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I632 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5118), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I633 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4441), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5071), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5118), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4441), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I636 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4414), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4237), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5071), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I637 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N489), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4858), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4414), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I638 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8830), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8675), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N489), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[27]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I639 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9231), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[28]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8830));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I640 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I641 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I642 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I643 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4591), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I644 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4623), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I645 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4765), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4591), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4623), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I646 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4440), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I647 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I648 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4544), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I649 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4394), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4440), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4544), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I650 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4412), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4765), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4394), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I651 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4937), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I652 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4635), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4937), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I653 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I654 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I655 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5152), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I656 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4812), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4635), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5152), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I657 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4446), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517), .A0(a_man[17]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5013), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4624), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4446), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5013), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I661 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4989), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4812), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4624), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N487), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4412), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4989), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4299), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4365), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4299), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I666 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4398), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I667 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4542), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4365), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4398), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I669 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4215), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I671 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I672 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4330), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4173), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4215), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4330), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4191), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4542), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4173), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I675 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4708), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I676 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4410), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4708), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I677 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4932), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4590), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4410), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4932), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I679 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4224), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I680 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I681 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4792), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I682 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4399), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4224), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4792), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4764), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4590), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4399), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N486), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4191), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4764), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I686 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4148), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I687 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4799), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I688 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4178), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4799), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4328), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4148), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4178), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I690 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I691 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4222), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I692 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5012), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4222), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I693 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5129), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I694 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4972), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5012), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5129), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I695 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4987), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4328), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4972), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I696 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4187), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I697 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5005), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I698 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4702), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5005), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I699 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4364), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4187), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4702), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I700 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I701 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5021), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I702 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4565), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4179), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5021), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4565), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I704 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4541), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4364), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4179), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I705 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N485), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4987), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4541), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I706 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4945), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I707 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4977), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I708 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5126), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4945), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4977), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I709 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4791), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I710 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I711 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I712 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4902), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I713 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4746), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4791), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4902), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I714 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4763), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5126), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4746), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I715 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4984), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4465), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4486), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4465), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I719 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4147), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4984), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4486), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I721 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4800), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I723 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I724 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4347), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I725 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4978), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4800), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4347), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I726 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4327), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4147), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4978), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I727 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N484), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4763), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4327), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I728 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I729 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4716), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I730 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4752), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I731 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4899), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4716), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4752), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I733 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4564), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I734 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5052), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I735 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4678), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5052), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I736 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4522), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4564), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4678), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I737 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4539), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4899), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4522), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I738 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I739 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4760), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I740 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I741 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4264), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I742 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4944), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4264), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4574), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4425), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I746 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4320), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I747 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5147), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4425), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4320), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I748 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4753), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4574), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5147), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I749 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5125), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4944), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4753), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I750 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N483), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4539), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5125), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I751 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4500), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I752 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4526), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I753 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4676), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4500), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4526), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I754 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5097), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I755 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4346), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5097), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I756 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4456), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I757 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4306), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4346), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4456), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I758 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4326), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4676), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4306), .B1(a_man[21]));
AO22XL float_div_cynw_cm_float_rcp_E8_M23_1_I759 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5007), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I760 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5007));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I762 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4537), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I763 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5040), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I764 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5058), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5040), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I765 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4715), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4537), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5058), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I766 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I767 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4353), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I768 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B(a_man[17]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I769 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I770 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4928), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I771 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4527), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4353), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4928), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I772 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4898), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4715), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4527), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I773 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N482), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4326), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4898), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I774 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I775 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4282), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I776 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I777 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4312), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I778 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4454), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4282), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4312), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I779 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5146), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I781 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4235), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I782 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5104), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5146), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4235), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I783 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5123), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4454), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5104), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I785 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4322), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I786 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4836), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I787 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4499), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4322), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4836), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4558), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I789 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I790 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5153), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4558), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I791 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4698), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I792 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4313), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5153), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4698), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I793 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4675), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4499), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4313), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I794 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N481), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5123), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4675), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I795 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4773), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I796 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5073), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4773), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4363), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I798 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5109), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4363), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I799 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4230), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5073), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5109), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I800 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4927), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I801 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I802 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5032), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I803 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4878), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4927), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5032), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I804 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4895), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4230), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4878), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I805 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5119), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I806 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I807 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4612), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I808 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4281), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5119), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4612), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I809 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4933), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I810 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4556), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I811 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4481), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4556), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I812 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5110), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4933), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4481), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I813 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4453), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4281), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5110), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I814 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N480), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4895), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4453), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I815 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4629), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I816 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4661), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I817 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4807), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4629), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4661), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I818 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4782), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I819 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4480), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4782), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I820 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4588), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I821 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4430), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4480), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4588), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I822 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4451), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4807), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4430), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I823 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4986), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4672), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4986), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I825 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4168), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I826 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4850), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4672), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4168), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I827 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4985), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I828 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4487), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4985), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I829 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5054), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4662), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4487), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5054), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I831 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5027), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4850), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4662), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I832 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4451), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5027), .B1(a_man[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I833 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I834 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4851), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I835 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I836 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4883), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I837 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5028), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4851), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4883), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I838 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I839 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4697), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I840 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4810), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I841 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4657), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4697), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4810), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I842 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4673), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5028), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4657), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I843 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4891), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I844 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4388), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I845 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5072), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4891), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4388), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I846 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I847 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4703), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I848 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4259), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4884), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4703), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4259), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I850 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4229), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5072), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4884), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I851 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N479), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4673), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4229), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I852 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8588), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26236), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N479));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I853 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9157), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8994), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N480), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8588));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I854 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8970), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8792), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N481), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9157));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I855 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8767), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8605), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N482), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8970));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I856 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8574), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9172), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N483), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8767));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I857 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9142), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8980), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N484), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8574));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I858 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8953), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8777), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N485), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9142));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I859 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8754), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8586), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N486), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8953));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I860 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8893), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8731), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N487), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8754));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I861 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I862 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4813), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I863 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4845), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I864 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4990), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4813), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4845), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I865 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4318), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I866 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4663), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4318), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I867 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I868 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4767), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I869 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4618), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4663), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4767), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I870 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4639), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4990), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4618), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I871 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4854), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I872 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4352), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I873 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5035), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4854), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4352), .B1(a_man[20]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I874 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4671), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I875 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I876 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4216), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I877 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4846), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4671), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4216), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I878 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4192), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5035), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4846), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I879 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N488), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4639), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4192), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I880 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7046), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I881 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4916), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I882 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4797), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4916), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I883 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4381), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I884 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4525), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4797), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4381), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I885 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I886 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4912), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I887 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4201), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4912), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I888 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5098), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I889 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4887), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5098), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I890 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4157), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4201), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4887), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I891 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4617), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4525), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4157), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I892 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I893 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4742), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I894 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4688), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I895 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4569), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4742), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4688));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I896 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4780), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I897 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4910), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I898 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4608), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4780), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4910));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I899 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4749), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4569), .B0(a_man[21]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4608));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I900 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[7]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4617), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .B0(a_man[22]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4749));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I901 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7271), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[7]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I902 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5075), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I903 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5018), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5075), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I904 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4607), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I905 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4750), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5018), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4607), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I906 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4420), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I907 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5113), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I908 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4375), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4420), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5113), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I909 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4839), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4750), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4375), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I910 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4966), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I911 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4913), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I912 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4796), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4966), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4913));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I913 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5002), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I914 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4190), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5137), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4190), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4831), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5002), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5137));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4974), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4796), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4831), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I918 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[8]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4839), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4974), .B1(a_man[22]));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I919 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[8]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I920 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7244), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I921 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7616), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7422), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7046), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7271), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7244));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I922 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7105), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I923 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7075), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I924 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7133), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I925 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7121), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6923), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7105), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7075), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7133));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I926 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7712), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7519), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7616), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6856), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7121));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I927 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7535), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7340), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7068), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7563), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7712));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I928 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7014), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I929 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6986), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I930 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .A(a_man[4]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I931 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7227), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7039), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7014), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6986), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I932 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7487), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I933 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7458), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_1_I934 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .A(a_man[3]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I935 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7023), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6834), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7487), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7458), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I936 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7518), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I937 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I938 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4570), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496), .B0(a_man[17]), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I939 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4163), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I940 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4311), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4570), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4163));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4996), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4665), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I943 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4956), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4996), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4665), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I944 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4393), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4311), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4956), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I945 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I946 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4518), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I947 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I948 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4466), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I949 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4351), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4518), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4466));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I950 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I951 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5060), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I952 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4554), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5060), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I953 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4686), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I954 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4383), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4554), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4686), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I955 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4524), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4351), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4383), .B1(a_man[21]));
AOI22X2 float_div_cynw_cm_float_rcp_E8_M23_1_I956 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[6]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4393), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4524), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I957 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6891), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I958 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6837), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I959 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7407), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7214), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7518), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6891), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6837));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I960 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7005), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7697), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7039), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7023), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7407));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I961 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7574), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I962 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7545), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I963 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7325), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7132), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7574), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7545), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I964 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7661), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I965 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7571), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I966 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7602), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I967 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7294), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7104), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7661), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7571), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7602));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I968 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I969 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6859), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I970 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7542), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I971 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I972 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7690), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I973 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6910), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7601), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6859), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7542), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7690));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I974 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7388), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7196), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7294), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6910), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7422));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I975 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7598), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7401), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7005), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7132), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7388));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7189), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7216), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7157), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I979 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7507), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7311), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7189), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7216), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7157));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I980 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7045), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5151), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I982 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I983 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4961), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I984 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5107), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5151), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4961), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I985 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4771), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I986 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4442), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I987 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4729), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4771), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4442), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4171), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5107), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4729), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I989 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4304), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I990 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4452), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I991 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4242), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4452), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I992 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5150), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4304), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4242));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I993 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4340), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I994 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4464), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I995 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4164), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4340), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4464), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I996 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4310), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5150), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4164), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I997 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[5]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4171), .B0(a_man[22]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4310));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I998 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7386), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[5]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I999 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7315), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7123), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7045), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7386));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1000 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7630), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1001 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7682), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7490), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7315), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7630), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6834));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1002 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6893), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7582), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7311), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6923), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7682));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1003 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7460), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1004 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7664), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[8]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1005 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7489), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1006 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7437), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7240), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7460), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7664), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7489));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1007 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7633), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1008 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7520), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1009 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7604), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1010 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6937), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7629), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7633), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7520), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7604));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1011 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7208), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7018), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7507), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7240), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7629));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1012 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7101), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6904), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6893), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7519), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7018));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1013 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7419), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7223), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7340), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7598), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7101));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1014 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7149), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6953), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6937), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7437), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7325));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1015 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7468), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7268), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7149), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7000), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7383));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1016 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7035), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6843), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7208), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7454), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6953));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1017 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6964), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7660), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6887), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7535), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7035));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1018 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[26]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7419), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7268), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7660));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1019 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9029), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8862), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8893), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N488), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[26]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1020 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[27]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6964), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7468), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7706));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1021 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9003), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9029), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[27]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8675));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1022 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1023 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1024 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8589), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1025 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9030), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8768), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1026 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4439), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1027 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4429), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4439), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634));
OR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1028 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4429));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I1029 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1030 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1031 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1032 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3661), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1033 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3683), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1034 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3421), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1035 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3661), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3683), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3421));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1036 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1037 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3629), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1039 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3546), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1040 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3750), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3676), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3664), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1043 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3743), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3663), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3750), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3676), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3664));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1044 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3418), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1045 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3414), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1046 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3716), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1047 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3558), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3470), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3418), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3414), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3716));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1048 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3501), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1049 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3648), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1050 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3620), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1051 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3454), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3758), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3501), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3648), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3620));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1052 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3487), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13732), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1054 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3690), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1055 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3626), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3542), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3487), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13732), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3690));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1056 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3410), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3715), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3558), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3758), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3542));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1057 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3774), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1058 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3529), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3444), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3454), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3774), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3626));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1059 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3663), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3410), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1060 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3596), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1061 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3569), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1062 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3537), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1063 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3474), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3397), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3596), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3569), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3537));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3453), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3467), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1066 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3649), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3564), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3453), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3743));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1067 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3529), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3397), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3564));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1068 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1069 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3672), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1070 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3544), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1071 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3422), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1072 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3656), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26349), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3672), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3544), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3422));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1073 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26325), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26348), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1077 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3458), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1078 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3498), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1079 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3646), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1080 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26352), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26338), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3458), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3498), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3646));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1081 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3437), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26315), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26325), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26348), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26352));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1082 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3502), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3425), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3470), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3656), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3437));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3601), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3450), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1085 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3634), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1086 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3556), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1087 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3630), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1088 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3482), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26322), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3634), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3556), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3630));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1089 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3725), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3640), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3601), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3450), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3482));
ADDFHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1090 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3502), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3725), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3715));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1091 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1092 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3625), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3765), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1095 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3554), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1096 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3597), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3510), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3625), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3765), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3554));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1097 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3510), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3474), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3649));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1098 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3637), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1099 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3518), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3713), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3548), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1102 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3550), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3461), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3518), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3713), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3548));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1103 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3597), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3637), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3461));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3724), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3692), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1109 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3724), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3692), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3550));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1110 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1111 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3687), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3706), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1117 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26340), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26327), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3687), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3706));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26335), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571));
NOR2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3722), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
NOR2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3591), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3473), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1122 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26307), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26354), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3722), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3591), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3473));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1123 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26318), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26363), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26340), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26335), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26307));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1124 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3604), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26341), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26349), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26322), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26318));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1125 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3604), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3640), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3425));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26312), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3468), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3682), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3553), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3535), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1132 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3666), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3581), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3553), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3535));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1133 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26333), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3433), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3468), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3682), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3666));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1134 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26344), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26330), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26338), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26312), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26333));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1135 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26344), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26315), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26341));
NAND2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3641), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3749), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1140 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3761), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3681), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3749));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3729), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3772), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3525), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1144 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3547), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3457), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3729), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3772), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3525));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1145 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3612), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3532), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3581), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3761), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3547));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3698), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3691), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3507), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1149 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26314), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3744), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3698), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3691), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3507));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1150 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26359), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3598), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26327), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26354), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26314));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1151 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3433), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3612), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3598));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1152 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26363), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26330));
NAND2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694));
NAND2X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3549), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3741), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3735), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3434), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1161 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3416), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1162 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26598), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26583), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3416));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1163 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3428), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26626), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3741), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3735), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26598));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3562), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3583), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1166 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3643), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26601), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3562), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3583));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1167 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3517), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1168 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3718), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3628), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3643), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3517), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3681));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1169 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3428), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3457), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3628));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1170 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3718), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3744), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3532));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1172 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489), .A1N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1173 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3395), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3568), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3577), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1176 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26621), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26608), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3395), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3568), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3577));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1177 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26601), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26621), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26626));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3621), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3402), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3633), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1181 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26603), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26593), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3402), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3633));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1182 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26583), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26608));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26636), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3441), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3460), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1186 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26610), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3441), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3460));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26585), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1188 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26615), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26610), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26585), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26593));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26627), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26606), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26587), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3623), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3615), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3452), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3685), .AN(a_man[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603));
ADDHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1196 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3451), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3452), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3685));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1197 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26637), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3623), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3615), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3451));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26637));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26615));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26619), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1201 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3570), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3668), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1203 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3511), .AN(a_man[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1204 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3668), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3511));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3617), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_1_I1207 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3555), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3624), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3617), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3555), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3404), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3526), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673), .A1N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3624), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3404));
OAI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26611), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3570), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3526), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26638), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1213 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26579), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26619), .A1N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26611), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26638));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26581), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26627), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26606), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26587), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26579));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1215 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26594), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1216 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3753), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26636), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26581), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1217 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3540), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3621), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3753), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3540));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3710), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3483), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1221 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3710), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3483));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694));
AOI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486));
AOI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392));
OAI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I1236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I1239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3618), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627));
OA21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3424), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3618));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3608), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3424));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I1242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3459), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3608));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3549), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3459));
MX2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3629), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3546), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3466), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3466));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6329), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4563), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4543), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4209), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4543), .B1(a_man[21]));
AO22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4563), .A1(a_man[22]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4209));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6264), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3403), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I1257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3403));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1258 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3680), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1259 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3704), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1260 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3582), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3704), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3762), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3582));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512));
NAND2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3766), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3675), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589));
OAI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430));
OAI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3442), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720));
AOI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1269 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3684), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3442));
OAI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I1270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3766), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3675), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3684));
MX2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1271 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3680), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3762), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1272 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6182), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1273 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4738), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1274 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1275 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4923), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4738), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1276 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4329), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5006), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4923), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4329), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4922), .A(a_man[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N456), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5006), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4922), .B1(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N456));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6385), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6451), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1283 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6459), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6383), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6182), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6385), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6451));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1284 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6329), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6264), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6459));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1285 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9081), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8925), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[24]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8586), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[24]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7331), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7130), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7269), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1289 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7200), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7009), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7331), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7130), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7269));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1290 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .A(a_man[0]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1291 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .A(a_man[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7515), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1293 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7217), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7028), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7515));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7073), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7103), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1296 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7700), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7510), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7217), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7073), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7103));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7156), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7302), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7241), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1300 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7587), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7391), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7156), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7302), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7241));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1301 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7181), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6987), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7200), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7700), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7587));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1302 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7185), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1303 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1304 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7359), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1305 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7212), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1306 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7091), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6896), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7185), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7359), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7212));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1307 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7566), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7372), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7214), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7091), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7601));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1308 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7274), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7087), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7697), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7181), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7566));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6918), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1310 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7568), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6857), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1312 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7108), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6913), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6918), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7568), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6857));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1314 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6971), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1315 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7540), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4931), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1318 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5016), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1319 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4732), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5016), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4882), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4931), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4732));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5121), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4548), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5121), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1323 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1324 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4217), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1325 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4509), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4548), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4217), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1326 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4970), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4882), .B0(a_man[21]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4509));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1327 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5099), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1328 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4595), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1329 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4930), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5099), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4595), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5026), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5139), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5026), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1333 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4241), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1334 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4962), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5139), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4241), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5106), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4930), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4962), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[4]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4970), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5106), .B1(a_man[22]));
CLKBUFX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[4]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7003), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1339 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7606), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7410), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6971), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7540), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7003));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1340 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7477), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7279), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7108), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7606), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7123));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6888), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7600), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6835), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1344 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7493), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7298), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6888), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7600), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6835));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1345 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6945), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1346 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7658), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1347 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6992), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7685), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7028), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6945), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7658));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1348 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6974), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7669), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7493), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6992), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7510));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1349 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7071), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6875), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7477), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7104), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6974));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1350 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7666), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7472), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7071), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7196), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7582));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1351 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7486), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7289), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7401), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7274), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7666));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1352 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[25]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6843), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7486), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7223));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1353 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9221), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9054), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9081), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8731), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[25]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1354 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9221), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[26]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8862));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9003));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7686), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7625), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7100), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4701), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4243), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4512), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4243), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4660), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4701), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4512), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4449), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4336), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4449), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5014), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4293), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4336), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5014), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4744), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4660), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4293), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4876), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4368), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1371 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4700), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4876), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4368));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1372 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4804), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1373 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4914), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4804), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967));
AOI22X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5039), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4733), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4914), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5039), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1377 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4881), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4700), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4733), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1378 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[3]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4744), .B0(a_man[22]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4881));
CLKBUFX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[3]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7505), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7038), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1382 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7621), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7428), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7100), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7505), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7038));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1383 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7376), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7184), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7686), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7625), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7621));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1384 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7360), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7166), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7009), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7376), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7391));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1385 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7456), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7259), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7360), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7490), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6987));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7183), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1387 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7153), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1388 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7356), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1389 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7011), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7703), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7183), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7153), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1390 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7127), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1391 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7445), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1392 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7384), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1393 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7513), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7317), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7127), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7445), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7384));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7328), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7414), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7238), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1397 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7394), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7202), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7328), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7414), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7238));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1398 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6878), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7570), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7011), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7513), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7394));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1399 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6861), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7553), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6878), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6896), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7279));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1400 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6955), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7648), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6861), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7372), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6875));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1401 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7162), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6968), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7087), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7456), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6955));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1402 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7162), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6904), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7289));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1403 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8664), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9244), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8925), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[24]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[24]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1404 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9054), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[25]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8664));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8983), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6305), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26412), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1409 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4515), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4547), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4694), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4515), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4547), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4720), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5055), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5128), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4720), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5055), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26419), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4694), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5128), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26399), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26412), .A1(a_man[22]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26419));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1417 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26399));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6511), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1421 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3427), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1422 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3594), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1423 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3506), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3594));
MX2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1424 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3427), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3506), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6371), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1426 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6355), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6281), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6305), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6511), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6371));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4301), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1428 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4335), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1429 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4476), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4301), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4335), .B1(a_man[20]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4503), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4834), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1432 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4901), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4503), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4834), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1433 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4559), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4476), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4901), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4247), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4871), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4247), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4908), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4254), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4871), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4908), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1438 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N454), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4559), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4254), .B1(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1439 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N454));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1440 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6295), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3644), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1443 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3560), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592));
MX2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1444 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3644), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3560), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1445 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6225), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1446 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6428), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1447 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6442), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6365), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6295), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6225), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6428));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1448 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6237), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1449 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6502), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6427), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6442), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6237), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6281));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1450 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6383), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6355), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6502));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1451 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9267), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9110), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[23]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8777), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[23]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_1_I1452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7475), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7211), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7299), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1456 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6900), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7589), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7475), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7211), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7299));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1457 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7263), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7074), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6900), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6913), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7410));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1458 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7565), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1459 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7596), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1460 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4485), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1461 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4295), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1462 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4434), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4485), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4295));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1463 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4227), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1464 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4949), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5136), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4227), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4949));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4793), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5085), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5136), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4793), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4521), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4434), .B0(a_man[21]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5085));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1469 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4520), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4654), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4520), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1471 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4150), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1472 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4484), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4654), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4150));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1473 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4743), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1474 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4689), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4743), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1475 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4779), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1476 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4815), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4779), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4513), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4689), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4815), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4659), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4484), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4513), .B1(a_man[21]));
AOI22X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[2]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4521), .B0(a_man[22]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4659));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7120), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[2]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1481 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7532), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7337), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7565), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7596), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7266), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7001), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7622), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1485 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7031), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1486 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7032), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6841), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7001), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7622), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7031));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1487 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7283), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7095), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7532), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7266), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7032));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1488 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7652), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7459), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7298), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7685), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7283));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1489 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7247), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7057), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7263), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7669), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7652));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1490 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1491 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7090), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6941), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6884), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1494 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6919), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7610), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6941), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7090), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6884));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1495 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6969), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1496 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7655), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1497 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6914), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1498 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7416), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7221), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6969), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7655), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6914));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1499 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7061), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1500 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7684), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1501 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6833), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1502 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7303), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7113), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7061), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7684), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6833));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1503 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7675), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7481), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6919), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7416), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7303));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1504 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7171), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6977), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7428), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7703), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7317));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1505 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7152), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6957), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7675), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7184), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7171));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1506 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7634), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7441), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7152), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7166), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7553));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1507 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7342), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7150), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7259), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7247), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7634));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1508 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7342), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7472), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6968));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1509 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8848), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8690), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[23]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[23]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9110));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1510 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9267), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9244), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8848));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4226), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4263), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4226), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5089), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4213), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4263), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5089), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5024), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1517 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4909), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5024), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1518 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4566), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1520 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4861), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4909), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4566), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4305), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4213), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4861), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1522 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4427), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1523 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4950), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1524 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4262), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4427), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4950), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1525 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4467), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1526 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4450), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1527 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4553), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1528 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4593), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4450), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4553), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1529 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4296), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4467), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4593), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1530 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4433), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4262), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4296), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1531 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[1]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4305), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4433), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1532 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7615), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1533 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7180), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1534 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7442), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1535 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7433), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7237), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7615), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7180), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7442));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1536 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6854), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1537 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7555), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7503), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7411), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1540 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6934), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7626), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7555), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7503), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7411));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1541 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7691), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7499), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7433), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6854), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6934));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1542 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7556), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7365), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7589), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7202), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7691));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1543 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7538), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7344), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7570), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7556), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1544 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7206), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[2]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7585), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1547 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7473), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1548 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7320), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7129), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7206), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7585), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7473));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1549 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7264), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7235), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7296), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1552 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7708), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7517), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7264), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7235), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7296));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1553 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7190), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6996), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7320), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7337), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1554 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7382), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1555 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7531), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7352), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1557 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7204), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7015), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7382), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7531), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7352));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1558 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7575), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7381), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6841), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7204), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7610));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1559 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7063), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6865), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7095), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7190), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7575));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1560 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7043), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6847), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7063), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7459), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6957));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1561 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7138), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6943), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7057), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7538), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7043));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1562 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7138), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7648), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7150));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1563 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8718), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9294), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8980), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[22]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1564 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6360), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1565 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6497), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1566 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6348), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1567 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1568 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096));
MXI2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26111), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1571 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26111));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6415), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1573 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5043), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4648), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5043), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1575 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4287), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1576 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4683), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4287), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1577 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26095), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4648), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4683), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1578 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5094), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1579 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5134), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1580 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4255), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5094), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5134), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1581 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4610), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1582 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4677), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4610), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1583 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26089), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4255), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4677), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1584 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26100), .A0(a_man[22]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26095), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26089), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1585 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26100));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6420), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1587 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6379), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6306), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6348), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6415), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6420));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1588 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6253), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6176), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6497), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6360), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6379));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1589 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6283), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6216), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6489), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1592 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6189), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6453), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6283), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6216), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6489));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1593 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6399), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6323), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6365), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6189), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1594 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6427), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6253), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6399));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1595 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9042), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8881), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[22]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1596 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8690), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8718), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9042));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1598 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778), .A(N12969), .B(N12863));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1600 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4371), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1601 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5057), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4371), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1602 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5149), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4865), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5149), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5009), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5057), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4865), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1605 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4579), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1606 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4685), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4579), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1607 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4348), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1608 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4642), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4685), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4348), .B1(a_man[20]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1609 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5103), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5009), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4642), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1610 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4208), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1611 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4723), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616), .B1(a_man[19]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1612 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5056), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4208), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4723));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1613 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4244), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1614 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4339), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736), .B0(a_man[17]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1615 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4366), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4339));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1616 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5090), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4244), .B0(a_man[20]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4366));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1617 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4212), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5056), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5090), .B1(a_man[21]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1618 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[0]), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5103), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .B0(a_man[22]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4212));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1619 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6954), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7327), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7681), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7058), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7170), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1626 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7225), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7036), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7681), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7058), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7170));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1627 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7593), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7398), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6954), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7327), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7225));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1628 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7079), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6883), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7113), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7221), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7593));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1629 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7446), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7250), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7079), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7481), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6977));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1630 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7029), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6852), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1632 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6880), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1633 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7614), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7421), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7029), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6852), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6880));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7711), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7086), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1636 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6997), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1637 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6845), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7536), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7711), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7086), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6997));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1638 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7117), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1639 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6966), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1640 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6940), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1641 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7118), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6921), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7117), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6966), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6940));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1642 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7098), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6903), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7614), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6845), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7118));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1643 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7485), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7287), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7129), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7237), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7517));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1644 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7465), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7265), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7499), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7098), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7485));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1645 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1646 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7199), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1647 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6912), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1648 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7551), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1649 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7349), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1650 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7243), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7055), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7551), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7349));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1651 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7504), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7308), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7199), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6912), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7243));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1652 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6982), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7677), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7015), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7626), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7504));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1653 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6962), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7657), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6996), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6982), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7381));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1654 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6946), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7639), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7465), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7365), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6962));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1655 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7424), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7229), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7344), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7446), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6946));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1656 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7424), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7441), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6943));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1657 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8913), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8745), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9172), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[21]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3491), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662));
XNOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3491), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I1661 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[17]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6457), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3696), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3394), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559));
MX2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1666 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3696), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3394), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1667 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6392), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6324), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1669 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6493), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6417), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6457), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6392), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6324));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6274), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1671 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1672 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4649), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4682), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4829), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4649), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4682), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1675 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4632), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1676 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4165), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1677 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4234), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4632), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4165), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4919), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4829), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4234), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1679 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4597), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1680 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1681 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4323), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1682 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4203), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4597), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4323), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4857), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4186), .A0(a_man[17]), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4240), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4857), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4186), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1686 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4605), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4203), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4240), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1687 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N451), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4919), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4605), .B1(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1688 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N451));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6330), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1690 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6260), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1691 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6465), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1692 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6299), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6228), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6330), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6260), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6465));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1693 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6468), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6394), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6493), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6274), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6299));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1694 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6191), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1695 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6245), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1696 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1697 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3439), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1698 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3523), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1699 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485));
MX2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1700 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3439), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3523), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1701 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6310), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1702 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6327), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6255), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6245), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6310));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4872), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1704 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4907), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1705 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5050), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4872), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4907), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1706 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4951), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1707 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4386), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4951), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1708 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4455), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4386), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1709 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5142), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5050), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4455), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1710 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4819), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1711 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4538), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B0(a_man[19]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1712 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4422), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4819), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4538), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1713 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5079), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1714 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4463), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5079), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1715 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4828), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4422), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4463), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N452), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5142), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4828), .B1(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6397), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1719 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6447), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6374), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6191), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6327), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6397));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6199), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1721 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6269), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6473), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1723 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6510), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6436), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6269), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6199), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6473));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1724 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6204), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1725 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6342), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1726 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6407), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1727 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6318), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6247), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6204), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6342), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6407));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1728 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6277), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6200), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6447), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6436), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6247));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1729 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6486), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6409), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6468), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6453), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6277));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1730 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6339), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6265), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6318), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6510), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6306));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1731 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6486), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6339), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6323));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7292), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1733 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7643), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1734 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7323), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1735 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7631), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7439), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7292), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7643), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7323));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1736 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7647), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1737 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7527), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1738 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7470), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1739 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7583), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1740 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7522), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7326), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7527), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7470), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7583));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1741 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7002), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7695), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7631), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7647), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7522));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1742 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7699), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7409), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7673), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1746 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7020), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6832), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7699), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7409), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7673));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1747 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7500), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1748 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7613), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1749 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7440), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1750 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7135), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6939), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7500), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7613), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7440));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1751 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7385), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7193), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7020), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7135), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7036));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1752 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7369), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7175), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7002), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7398), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7385));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1753 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6889), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7580), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7421), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7536), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6921));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1754 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6870), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7561), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6903), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6889), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7287));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1755 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7348), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7155), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7369), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6883), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6870));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1756 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7333), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7142), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6865), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7250), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7348));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1757 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7333), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6847), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7229));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1758 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9098), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8942), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8605), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[20]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[20]));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1759 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9235), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9070), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[21]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9098));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1760 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8913), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9235), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8881));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1762 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4423), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1763 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4462), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1764 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4606), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4423), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4462), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1765 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4407), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1766 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4963), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1767 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5031), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4407), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4963), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1768 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4690), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4606), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5031), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1769 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4370), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1770 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5120), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1771 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5000), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4370), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5120), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1772 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4637), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1773 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4983), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1774 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5037), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4637), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4983), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1775 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4379), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5000), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5037), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1776 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N450), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4690), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4379), .B1(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1777 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N450));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1778 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6452), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1779 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6251), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6316), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1781 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6285), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6209), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6452), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6251), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6316));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1782 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6449), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1783 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6178), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6381), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1785 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6474), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6401), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6449), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6178), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6381));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1786 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6259), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6185), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6285), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6474), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6417));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1787 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6183), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6367), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1789 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6435), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1790 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6301), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1791 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6499), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6423), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6435), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6367), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6301));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1792 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6431), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6357), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6255), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6183), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6499));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1793 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6405), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6333), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6431), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6228), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6374));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1794 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6422), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6350), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6394), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6259), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6405));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1795 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6422), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6265), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6409));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1796 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7143), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6936), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1798 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7040), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6846), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7143), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6936));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1799 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7379), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1800 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7404), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7210), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7040), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7379), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7055));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1801 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7056), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1802 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7083), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1803 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6995), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1804 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6925), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7617), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7056), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7083), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6995));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1805 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7224), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1806 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7197), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1807 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7026), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1808 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7423), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7228), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7224), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7197), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7026));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1809 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7167), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1810 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7114), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1811 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6909), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1812 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7313), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7122), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7114), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6909), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7167));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1813 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6907), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7599), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6925), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7423), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7313));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1814 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7270), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7084), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7308), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7404), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6907));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1815 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7256), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7066), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7677), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7270), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7175));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1816 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6850), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7541), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7657), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7265), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7256));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1817 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6850), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7639), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7142));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1818 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9282), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9128), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8792), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[19]));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1819 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8680), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9257), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[20]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9282));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1820 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8680), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8745), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9070));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1821 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209));
CLKAND2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1822 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568), .A(N13035), .B(N12722));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1823 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26710), .A(N12754), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1825 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6373), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1826 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4204), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1827 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4239), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1828 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4380), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4204), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4239), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1829 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4185), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4735), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1831 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4809), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4185), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4735), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1832 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4472), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4380), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4809), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1833 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4153), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1834 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4892), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1835 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4776), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4153), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4892), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1836 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4189), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1837 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4758), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1838 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4814), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4189), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4758), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1839 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4161), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4776), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4814), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1840 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N449), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4472), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4161), .B1(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1841 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N449));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1842 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6239), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1843 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6440), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1844 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6455), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6380), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6373), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6239), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6440));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1845 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3763), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695));
CLKXOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1846 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3763));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1847 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6501), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1848 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6508), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6234), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1850 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6308), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6233), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6501), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6508), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6234));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1851 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6238), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6505), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6455), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6308), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6401));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1852 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6307), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1853 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1854 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3575), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1855 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3659), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508));
MX2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1856 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3575), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3659), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1857 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6353), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1858 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6424), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1859 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6220), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1860 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6336), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6262), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6353), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6424), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6220));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1861 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6494), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1862 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26090), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1863 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26108), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104));
NOR3X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1864 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6358), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26090), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26108));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1865 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6287), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1866 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6482), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6408), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6494), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6358), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6287));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1867 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6267), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6190), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6307), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6336), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6482));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1868 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6386), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26219), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6267), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6209), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6357));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1869 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6214), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6480), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6238), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6185), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6386));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1870 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6214), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6200), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6350));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1871 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7255), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1872 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7282), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1873 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6963), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1874 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7698), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7508), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7255), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7282), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6963));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1875 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7291), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7102), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7439), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7698), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7326));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1876 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7662), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7469), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7695), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7291), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7193));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1877 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7611), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1878 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7406), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1879 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7215), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7025), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7406));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1880 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7526), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1881 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7550), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1882 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7467), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1883 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7106), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6911), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7526), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7550), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7467));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1884 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7198), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7006), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6846), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7215), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7106));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1885 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7679), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7488), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6832), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6939), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7198));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1886 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7640), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1887 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7581), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1888 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6869), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1889 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7491), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7295), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7640), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7581), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6869));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1890 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7670), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1891 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7696), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1892 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7495), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1893 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7603), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7408), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7670), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7696), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7495));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1894 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7584), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7389), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7491), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7603), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7228));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1895 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6844), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1896 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7436), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1897 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7194), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1898 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7052), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1899 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6899), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7588), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7194), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7052));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1900 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6989), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7683), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6844), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7436), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6899));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1901 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7088), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6894), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7122), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7617), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6989));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1902 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7178), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6985), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7584), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7210), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7088));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1903 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7158), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6965), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7580), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7679), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7178));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1904 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7644), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7452), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7561), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7662), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7158));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1905 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26263), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7644), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7155), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7541));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1906 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8733), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9307), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8994), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[18]));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1907 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8866), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8707), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[19]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8733));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1908 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8866), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8942), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9257));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1909 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1910 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6498), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1911 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6291), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1912 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6430), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1913 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6289), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6217), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6498), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6291), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6430));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1914 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6413), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6341), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6289), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6423), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6233));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6226), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6344), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6278), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1918 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6507), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6432), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6344), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6278));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I1919 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1920 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1921 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6206), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1922 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6478), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1923 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6211), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1924 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6315), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6242), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6206), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6478), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6211));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1925 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6438), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6361), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6226), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6507), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6315));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1926 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6411), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1927 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6416), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1928 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6484), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1929 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6464), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6389), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6411), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6416), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6484));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1930 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6349), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1931 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6403), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1932 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6470), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1933 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6490), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6414), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6470), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1934 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6284), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1935 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6273), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6196), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6349), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6284), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6490));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1936 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6249), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6512), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6464), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6273), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6262));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1937 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6223), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6488), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6438), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6380), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6249));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1938 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26266), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26253), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6505), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6413), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6223));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1939 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26243), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26266), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6333), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6480));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1940 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7251), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7277), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7081), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1943 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7281), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7093), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7251), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7277), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7081));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1944 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7111), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1945 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7141), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1946 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7222), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1947 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7672), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7479), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7111), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7141), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7222));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1948 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7374), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7182), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7281), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7025), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7672));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1949 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7474), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7275), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7374), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7508), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7006));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1950 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7564), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7371), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7599), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7102), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7474));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1951 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7546), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7353), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7084), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7564), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7469));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1952 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26250), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26233), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7546), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7066), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7452));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1953 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8928), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26198), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26250), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26236), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26263));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1954 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9056), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8898), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8928), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[18]));
ADDFHXL float_div_cynw_cm_float_rcp_E8_M23_1_I1955 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9056), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9128), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8707));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1956 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833));
CLKAND2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I1957 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092), .A(N12983), .B(N12737));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1958 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7341), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1959 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7165), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1960 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7312), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1961 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7169), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6975), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7341), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7165), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7312));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1962 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6876), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7567), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7408), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7169), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6911));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1963 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7668), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1964 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7524), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1965 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6960), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7654), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7668), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7524));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1966 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7021), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1967 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7554), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7362), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6960), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7021), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7588));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1968 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7260), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7072), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7554), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7295), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7683));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1969 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6970), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7667), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7389), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6876), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7260));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I1970 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7069), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6873), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6970), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7488), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6985));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1971 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26216), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26203), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7069), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6965), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7353));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I1972 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8840), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1973 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1974 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4403), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1975 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4436), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4583), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4403), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4436), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4258), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4362), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1979 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4210), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4258), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4362), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1980 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4228), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4583), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4210), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4447), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1982 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4965), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1983 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4628), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4447), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4965), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1984 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4761), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1985 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4265), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4761), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1986 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4833), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1987 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4437), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4265), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4833), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4806), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4628), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4437), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I1989 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N477), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4228), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4806), .B1(a_man[22]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I1990 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7694), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1991 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7608), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1992 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7578), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1993 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6848), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7539), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7694), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7608), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1994 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6842), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1995 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6866), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1996 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7548), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I1997 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7346), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7154), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6866), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7548), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6842));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1998 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6924), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I1999 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7637), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2000 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6897), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2001 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7232), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7044), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6924), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7637), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2002 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7060), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6863), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6848), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7346), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7232));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2003 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7444), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7248), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7479), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7093), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6975));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2004 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7650), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7457), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7182), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7060), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7444));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2005 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7357), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7164), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7650), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6894), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7275));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2006 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[15]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[14]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7371), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7357), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6873));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2007 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26240), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26222), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N477), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[15]));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2008 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26230), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26214), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26216), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8840), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26240));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2009 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6332), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2010 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6266), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2011 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6337), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2012 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6296), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6224), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6332), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6266), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6337));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2013 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6195), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2014 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6201), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2015 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6270), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2016 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6444), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6370), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6195), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6201), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6270));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2017 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6419), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6345), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6432), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6296), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6444));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2018 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6396), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6319), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6217), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6408), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6419));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2019 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26246), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26229), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6190), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6396), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6341));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2020 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26225), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26211), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26246), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26219), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26253));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2021 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9246), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26227), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26230), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26225), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26243));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2022 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9246), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9307), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8898));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2023 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2024 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6475), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2025 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6257), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2026 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6188), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2027 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6279), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6203), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6257), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2028 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6256), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6181), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6475), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6279), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6414));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2029 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6230), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6496), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6256), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6242), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6389));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2030 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6202), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6469), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6230), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6361), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6512));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2031 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26206), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[15]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6488), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6202), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26229));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2032 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26260), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26247), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26214), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26233), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26206));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2033 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26260), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26198), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26227));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2034 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223));
CLKAND2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2035 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859), .A(N12742), .B(N12990));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2036 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2037 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6393), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6320), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2039 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6326), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2040 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6235), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6500), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6393), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6320), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6326));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6454), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6387), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2043 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6458), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2044 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6425), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6351), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6454), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6387), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6458));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2045 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6402), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6328), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6235), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6425), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6224));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2046 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6376), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6302), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6402), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6196), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6345));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2047 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26213), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[14]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6376), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6319), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6469));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2048 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7249), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2049 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7276), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2050 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7413), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7220), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7249), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7276));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2051 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7309), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2052 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7338), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7137), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2054 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6916), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7607), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7309), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7338), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7137));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2055 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7620), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7427), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7654), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7413), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6916));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2056 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7161), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2057 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7191), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2058 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7219), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2059 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7300), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7110), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7161), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7191), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2060 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7125), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6927), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7539), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7300), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7154));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2061 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6944), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7636), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7362), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7620), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7125));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2062 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7151), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6956), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6944), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7567), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7072));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2063 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[13]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7667), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7151), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7164));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7366), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7392), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2066 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6839), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2067 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6864), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2068 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7367), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7173), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6839), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6864));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2069 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7689), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7497), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7366), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7392), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2070 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6895), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2071 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6922), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2072 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7692), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2073 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6868), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7559), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6922), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7692), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6895));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7632), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7665), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6978), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2077 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7253), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7064), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7632), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7665), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6978));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2078 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7187), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6994), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7220), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6868), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7253));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2079 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7512), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7316), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7044), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7689), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7187));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2080 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7330), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7140), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7512), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6863), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7248));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2081 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[12]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7457), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7330), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6956));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2082 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6179), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6445), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6437), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2085 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6503), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2086 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6304), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6231), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6437), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6503));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2087 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6174), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26496), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6179), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6445), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6304));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2088 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6192), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6456), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6351), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6174), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6500));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2089 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6378), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2090 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6311), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2091 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6218), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6483), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6378), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6311));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2092 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26415), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26417), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_1_I2094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6241), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26415), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26417));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2095 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6513), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2096 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6246), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2097 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6363), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6290), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6241), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6513), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6246));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2098 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6382), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6309), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6203), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6218), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6363));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2099 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6210), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6476), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6382), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6370), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6181));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2100 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[12]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6328), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6192), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6476));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2101 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8747), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8575), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[13]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[13]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2102 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[13]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6210), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6302));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2103 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8657), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9236), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[14]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[14]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[14]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2104 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[14]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8747), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9236));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2105 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26200), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8720), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26203), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26222), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26213));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2106 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8657), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8720));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I7811 (.Y(N13125), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I7812 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26563), .A(N13132));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6951), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2109 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7306), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2110 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7335), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2111 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7705), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7514), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7306), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7335));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2112 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7641), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7449), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6951), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7705), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7173));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2113 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7572), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7378), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7110), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7607), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7641));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2114 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7010), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7702), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7572), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7427), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6927));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2115 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[11]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7636), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7010), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7140));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6362), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6297), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6369), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2119 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26489), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26473), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6362), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6297), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6369));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2120 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6321), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26455), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26489), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6483), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6290));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2121 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[11]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6309), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6321), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6456));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2122 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8835), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8683), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[12]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[12]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[12]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2123 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[13]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8835), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8575));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26548), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7453), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7245), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7420), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2128 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7590), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7396), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7453), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7245), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7420));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7363), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7390), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7272), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2132 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7203), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7012), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7363), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7390), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7272));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2133 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7145), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6949), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7590), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7203), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7559));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2134 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7077), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6881), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7145), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7497), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6994));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2135 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26468), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7316), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7077), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7702));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6892), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6920), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2138 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7543), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7351), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6892), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6920));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6948), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6976), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6860), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2142 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7047), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6851), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6948), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6976), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6860));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2143 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7096), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6901), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7514), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7543), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7047));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2144 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7529), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7334), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7096), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7064), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7449));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2145 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26452), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26439), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7378), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7529), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6881));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6491), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6421), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6354), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2149 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26499), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26483), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6491), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6421), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6232), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6288), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6222), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2153 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6197), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6466), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6288), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6222));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2154 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26449), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26504), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6197), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6232), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6231));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2155 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26479), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26464), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26473), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26499), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26504));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2156 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9035), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26481), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26452), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26479), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26468));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2157 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8946), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8770), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[11]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[11]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9035));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2158 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[12]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8946), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8683));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8769), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2160 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26486), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26496), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26449), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26455));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2161 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[11]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[11]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8770));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2162 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9199), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7418), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7450), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7509), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2166 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7267), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7080), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7418), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7450), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7509));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2167 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6931), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7623), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7351), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7267), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6851));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2168 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7007), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2169 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7037), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2170 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7358), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7387), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2172 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6886), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7577), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7358), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7387));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2173 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7430), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7234), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7007), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7037), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6886));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2174 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7483), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7284), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7430), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7012), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7396));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2175 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26461), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6931), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6901), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7284));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6412), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6275), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2178 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6243), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6412), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6275));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7034), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6972), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2181 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7501), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7305), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7034), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6972));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7480), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2183 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7659), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7466), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7501), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7480), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7577));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2184 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[7]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7234), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7659), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7623));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7094), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7004), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7065), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2188 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6999), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7094), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7004), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7065));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2189 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[6]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7080), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6999), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7466));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2193 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8760), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[5]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2194 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8671), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[6]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8760));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2195 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26444), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[7]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8671));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2196 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26474), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26483), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26461), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6479), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6207), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6334), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6268), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2201 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6433), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6334), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6268));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2202 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6390), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6479), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6207), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6433));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2203 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26458), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6243), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6466), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6390));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2204 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26493), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6949), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7483), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7334));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2205 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26436), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26490), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26458), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26493), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26439));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2206 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26464), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26474), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26490));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2207 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8607), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26436), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26481), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26486));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9283), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2210 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9190), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7506), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7476), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2213 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7612), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7417), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7506), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7476));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7534), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2215 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7558), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2216 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7115), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7534), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7558), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7417));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2217 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[5]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7305), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7612), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7115));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2218 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9088), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9190), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[5]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[5]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2219 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8999), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[6]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9088));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2220 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8901), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[7]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8999));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2221 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[8]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[8]), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8901));
AND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8971), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9059), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8734), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9158), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8822), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7089), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7148), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2229 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[3]), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7089), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7148));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9248), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8931), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[2]));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8655), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885), .C(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310), .D(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8756), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[2]));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9210), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8931), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8655), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8756));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8926), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9248), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9210), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[3]), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8668), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8636), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8822), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8926), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8668));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9006), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9158), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8636), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8562), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8617), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8734), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9006), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8562));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8892), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9059), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8617), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8639), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9165), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061), .A1N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8892), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8639));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8795), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8579), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8971), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9165), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8795));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9130), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8762), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9283), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8579), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9130));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8868), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8607), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8708), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8607), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8836), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8762), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8868), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8708));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9034), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8930), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9199), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8836), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9034));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8606), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26553), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8769), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8930), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8606));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8944), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807));
AOI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I2257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26561), .A0(N13070), .A1(N13072), .B0(N13068));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2258 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26565), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562));
OAI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I2259 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26563), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26561), .B0(N13013));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_1_I2260 (.CO(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019), .S(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26200), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26211), .CI(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26247));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8873), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667));
AND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632), .A(N13023), .B(N12687));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8715), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9038), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9288), .A0(N12682), .A1(N13023), .B0(N13146));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9288));
AOI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I2268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2269 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8949), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2271 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9202), .A0(N12744), .A1(N12990), .B0(N13142));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2272 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9202));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2273 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2274 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8839), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2275 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13738), .A0(N12983), .A1(N12739), .B0(N13138));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2276 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13738));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598));
OAI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I2278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053));
NOR2X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179), .A(N13106), .B(N13108));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8750), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9010), .A0(N13035), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179), .B0(N13134));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_1_I2282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9010));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9003));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8806), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2289 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622), .A0(N12969), .A1(N12719), .B0(N12967));
AOI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I2290 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2291 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2293 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9185), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8589), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9185));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2300 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2302 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2303 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8793), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2304 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8604), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8793));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2305 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8861), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8768), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8604));
OAI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26703), .A0(N13644), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964), .B0(N12752));
AOI21X4 float_div_cynw_cm_float_rcp_E8_M23_1_I2307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26710), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26703));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[39]), .A(N12500), .B(N12502), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2309 (.Y(x[22]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[39]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2310 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8601), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9242), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8601));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9080), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2314 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[38]), .A(N12493), .B(N12495), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2315 (.Y(x[21]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[38]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8752), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2318 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8584), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2319 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[37]), .A(N12486), .B(N12488), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2320 (.Y(x[20]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[37]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I2322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2323 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8736), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2324 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8736), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2325 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8665), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2326 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9015), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8665));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2327 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8846), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2328 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165), .A(N12896), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2329 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2333 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122));
OAI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2334 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156), .A0(N12896), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622), .B0(N12894));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26140), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26140));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[35]), .A(N12479), .B(N12481), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2340 (.Y(x[18]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[35]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9112), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9265), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9112));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9108), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2345 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[34]), .A(N12472), .B(N12474), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2346 (.Y(x[17]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[34]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2347 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2348 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8774), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2349 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8616), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2350 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[33]), .A(N12465), .B(N12467), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2351 (.Y(x[16]), .A0(N13648), .A1(N13650), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[33]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I2353 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26737), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2354 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26143), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26168), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26143));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26149), .A0N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151), .A1N(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26168));
MXI2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[32]), .A(N12549), .B(N12547), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26149));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2358 (.Y(x[15]), .A0(N13648), .A1(N13650), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[32]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8746), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I2360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9086), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9086), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9174), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9040), .A(N12747), .B(N12749));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8879), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8746), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8743), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8570), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8743), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8570));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9040), .B(N12544), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2371 (.Y(x[14]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[31]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2372 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9198), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2373 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8867), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9292), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8867));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9140), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9198), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[30]), .A(N12535), .B(N12537), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2377 (.Y(x[13]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[30]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2378 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9008), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8803), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9008), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8651), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9008), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[29]), .A(N12528), .B(N12530), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2382 (.Y(x[12]), .A0(N13648), .A1(N13650), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[29]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9259), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2384 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[28]), .A(N12574), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2385 (.Y(x[11]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[28]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9247), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I2387 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9065), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2388 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8696), .A(N12834), .B(N12719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2389 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8696), .B(N12942));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_1_I2390 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8929), .A0(N12834), .A1(N12863), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2391 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9068), .A(N13456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8929));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2392 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8911), .A(N13456), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011));
INVXL float_div_cynw_cm_float_rcp_E8_M23_1_I2393 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9167), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9004), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635));
AOI21X2 float_div_cynw_cm_float_rcp_E8_M23_1_I2396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612), .A0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903), .A1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9167), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9004));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9068), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8911), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2398 (.Y(x[10]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[27]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8956), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8625), .A(N12863), .B(N12719));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8572), .A(N12712), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8625));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9170), .A(N12712), .B(N12719));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8572), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9170), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2404 (.Y(x[9]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[26]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9284), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8831), .A(N13460), .B(N12729));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8677), .A(N13460), .B(N12734));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8831), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8677), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2409 (.Y(x[8]), .A0(N13650), .A1(N13648), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[25]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8796), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[24]), .A(N12554), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2412 (.Y(x[7]), .A0(N13648), .A1(N13650), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[24]));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060), .AN(N13134), .B(N13035));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8940), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9096), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060), .B(N12722));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8940), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9096), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2417 (.Y(x[6]), .A0(N13648), .A1(N13650), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[23]), .B1(N13646));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8563), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179), .B(N12722));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8563));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2420 (.Y(x[5]), .A0(N13648), .A1(N13650), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[22]), .B1(N13646));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2421 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823), .AN(N13138), .B(N12983));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2422 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9195), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823), .B(N12739));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2423 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8602), .A(N12737), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2424 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9195), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8602), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2425 (.Y(x[4]), .A0(N13648), .A1(N13650), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[21]), .B1(N13646));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9087), .AN(N12739), .B(N12737));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9087));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2428 (.Y(x[3]), .A0(N13648), .A1(N13650), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[20]), .B1(N13646));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2429 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592), .AN(N13142), .B(N12990));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8705), .A(N12744), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8863), .A(N12742), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2432 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13851), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2433 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13851));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8705), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8863), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2435 (.Y(x[2]), .A0(N13648), .A1(N13650), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[19]), .B1(N13646));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8854), .AN(N12744), .B(N12742));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8854), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2438 (.Y(x[1]), .A0(N13648), .A1(N13650), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[18]), .B1(N13646));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2439 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117), .AN(N13146), .B(N13023));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2440 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8967), .A(N12682), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_1_I2441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9126), .A(N12687), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8967), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9126), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2443 (.Y(x[0]), .A0(N13648), .A1(N13650), .B0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[17]), .B1(N13646));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_1_I2444 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26692), .AN(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2445 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26698), .A(N12569), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_1_I2446 (.Y(x[19]), .A0(N13648), .A1(N13650), .B0(N13646), .B1(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26698));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2447 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2448 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2449 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[7]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2450 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[6]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[5]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[4]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[3]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[2]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[1]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_1_I2456 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[0]), .S0(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_1_I2457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[31]), .AN(a_sign), .B(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29));
reg x_reg_23__I2481_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__I2481_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[23];
	end
assign x[23] = x_reg_23__I2481_QOUT;
reg x_reg_24__I2482_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__I2482_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[24];
	end
assign x[24] = x_reg_24__I2482_QOUT;
reg x_reg_25__I2483_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_25__I2483_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[25];
	end
assign x[25] = x_reg_25__I2483_QOUT;
reg x_reg_26__I2484_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__I2484_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[26];
	end
assign x[26] = x_reg_26__I2484_QOUT;
reg x_reg_27__I2485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__I2485_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[27];
	end
assign x[27] = x_reg_27__I2485_QOUT;
reg x_reg_28__I2486_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__I2486_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[28];
	end
assign x[28] = x_reg_28__I2486_QOUT;
reg x_reg_29__I2487_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__I2487_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[29];
	end
assign x[29] = x_reg_29__I2487_QOUT;
reg x_reg_30__I2488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I2488_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[30];
	end
assign x[30] = x_reg_30__I2488_QOUT;
reg x_reg_31__I2489_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I2489_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[31];
	end
assign x[31] = x_reg_31__I2489_QOUT;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[0] = x[0];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[1] = x[1];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[2] = x[2];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[3] = x[3];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[4] = x[4];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[5] = x[5];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[6] = x[6];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[7] = x[7];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[8] = x[8];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[9] = x[9];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[10] = x[10];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[11] = x[11];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[12] = x[12];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[13] = x[13];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[14] = x[14];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[15] = x[15];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[19] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[20] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[21] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[22] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[23] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[24] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[36] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  srjwTQrdrho= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



