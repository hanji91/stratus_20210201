/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:37:56 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_3_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__9,
	inst_cellmath__10,
	inst_cellmath__11,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__16,
	inst_cellmath__17,
	inst_cellmath__18;
wire [8:0] inst_cellmath__27;
wire [7:0] inst_cellmath__29;
wire  inst_cellmath__30,
	inst_cellmath__31,
	inst_cellmath__32;
wire [49:0] inst_cellmath__33;
wire  inst_cellmath__34;
wire [7:0] inst_cellmath__35;
wire [49:0] inst_cellmath__36,
	inst_cellmath__37;
wire [25:0] inst_cellmath__39;
wire  inst_cellmath__42,
	inst_cellmath__43,
	inst_cellmath__44;
wire [26:0] inst_cellmath__45;
wire  inst_cellmath__48;
wire [5:0] inst_cellmath__49;
wire [24:0] inst_cellmath__50;
wire  inst_cellmath__54,
	inst_cellmath__55;
wire [23:0] inst_cellmath__57;
wire [9:0] inst_cellmath__59;
wire  inst_cellmath__62,
	inst_cellmath__63;
wire [22:0] inst_cellmath__64;
wire  inst_cellmath__66;
wire [7:0] inst_cellmath__68;
wire  inst_cellmath__70,
	inst_cellmath__71;
wire N547,N556,N557,N558,N559,N560,N561 
	,N562,N563,N565,N566,N567,N568,N569,N570 
	,N571,N572,N574,N575,N626,N627,N628,N630 
	,N631,N632,N633,N634,N635,N638,N642,N645 
	,N650,N651,N652,N653,N655,N658,N661,N662 
	,N663,N664,N665,N666,N667,N668,N669,N670 
	,N671,N672,N673,N674,N675,N676,N677,N706 
	,N710,N3083,N3085,N3106,N3114,N3117,N3119,N3123 
	,N3125,N3128,N3134,N3138,N3168,N3170,N3191,N3199 
	,N3202,N3204,N3208,N3210,N3213,N3219,N3223,N3269 
	,N3273,N3291,N3295,N3319,N3321,N3324,N3327,N3331 
	,N3333,N3338,N3343,N3348,N3352,N3358,N3364,N3367 
	,N3403,N3404,N3405,N3406,N3408,N3410,N3412,N3413 
	,N3414,N3415,N3416,N3419,N3420,N3421,N3423,N3424 
	,N3426,N3428,N3430,N3431,N3432,N3433,N3434,N3436 
	,N3437,N3439,N3441,N3443,N3444,N3446,N3447,N3449 
	,N3451,N3453,N3454,N3455,N3457,N3459,N3460,N3461 
	,N3462,N3465,N3467,N3468,N3470,N3471,N3473,N3475 
	,N3477,N3478,N3479,N3480,N3482,N3483,N3485,N3487 
	,N3488,N3489,N3490,N3492,N3494,N3495,N3496,N3498 
	,N3499,N3501,N3502,N3503,N3504,N3505,N3506,N3507 
	,N3508,N3511,N3512,N3513,N3515,N3517,N3518,N3520 
	,N3522,N3524,N3525,N3527,N3528,N3530,N3532,N3534 
	,N3535,N3536,N3537,N3539,N3540,N3541,N3542,N3544 
	,N3546,N3547,N3548,N3550,N3551,N3671,N3678,N3682 
	,N3686,N3688,N3691,N3694,N3698,N3701,N3729,N3730 
	,N3769,N3840,N3842,N3843,N3844,N3846,N3848,N3849 
	,N3851,N3852,N3853,N3855,N3857,N3858,N3859,N3860 
	,N3862,N3864,N3866,N3867,N3868,N3869,N3872,N3874 
	,N3876,N3877,N3879,N3881,N3883,N3884,N3885,N3886 
	,N3889,N3890,N3891,N3892,N3893,N3895,N3896,N3897 
	,N3899,N3901,N3902,N3904,N3906,N3907,N3909,N3911 
	,N3913,N3914,N3915,N3916,N3919,N3920,N3921,N3923 
	,N3925,N3926,N3927,N3928,N3930,N3932,N3934,N3935 
	,N3937,N3939,N3940,N3942,N3945,N3947,N3949,N3950 
	,N3951,N3952,N3954,N3956,N3958,N3959,N3960,N3962 
	,N3964,N3965,N3966,N3968,N3970,N3971,N3973,N3975 
	,N3977,N3978,N3979,N3980,N3983,N3984,N3985,N3986 
	,N3988,N3990,N3992,N3993,N3994,N3996,N3998,N3999 
	,N4001,N4003,N4005,N4006,N4007,N4008,N4011,N4012 
	,N4014,N4016,N4017,N4018,N4019,N4021,N4022,N4024 
	,N4026,N4027,N4029,N4031,N4032,N4033,N4034,N4035 
	,N4037,N4040,N4041,N4042,N4044,N4046,N4047,N4048 
	,N4049,N4051,N4053,N4055,N4056,N4277,N4332,N4333 
	,N4335,N4337,N4339,N4342,N4343,N4346,N4349,N4351 
	,N4353,N4354,N4356,N4362,N4363,N4366,N4371,N4372 
	,N4400,N4578,N4579,N4582,N4583,N4585,N4586,N4589 
	,N4593,N4594,N4595,N4597,N4600,N4603,N4604,N4609 
	,N4610,N4612,N4616,N4618,N4620,N4621,N4624,N4626 
	,N4628,N4635,N4636,N4639,N4643,N4644,N4647,N4648 
	,N4653,N4654,N4657,N4659,N4663,N4664,N4665,N4666 
	,N4667,N4668,N4672,N4673,N4676,N4677,N4679,N4682 
	,N4684,N4687,N4691,N4692,N4695,N4699,N4700,N4701 
	,N4704,N4706,N4707,N4709,N4713,N4717,N4718,N4719 
	,N4722,N4723,N4824,N4826,N4827,N4828,N4829,N4831 
	,N4832,N4835,N4836,N4837,N4838,N4840,N4841,N4842 
	,N4845,N4846,N4847,N4848,N4850,N4852,N4855,N4856 
	,N4857,N4859,N4860,N4862,N4863,N4864,N4866,N4868 
	,N4869,N4870,N4872,N4873,N4874,N4877,N4878,N4880 
	,N4881,N4883,N4885,N4887,N4888,N4889,N4891,N4892 
	,N4893,N4894,N4896,N4898,N4900,N4901,N4902,N4904 
	,N4905,N4907,N4909,N4910,N4911,N4913,N4914,N4917 
	,N4918,N5043,N5064,N5113,N5116,N5122,N5128,N5129 
	,N5131,N5132,N5134,N5135,N5137,N5138,N5139,N5141 
	,N5142,N5143,N5145,N5146,N5148,N5149,N5152,N5155 
	,N5157,N5159,N5161,N5162,N5164,N5165,N5166,N5168 
	,N5169,N5171,N5172,N5174,N5175,N5177,N5178,N5180 
	,N5181,N5183,N5186,N5189,N5191,N5192,N5193,N5195 
	,N5196,N5198,N5199,N5202,N5204,N5205,N5206,N5208 
	,N5210,N5211,N5213,N5214,N5216,N5217,N5218,N5220 
	,N5223,N5226,N5228,N5229,N5231,N5233,N5235,N5236 
	,N5238,N5239,N5240,N5242,N5243,N5245,N5247,N5248 
	,N5251,N5253,N5254,N5257,N5258,N5261,N5263,N5265 
	,N5266,N5267,N5269,N5270,N5272,N5274,N5275,N5278 
	,N5279,N5283,N5284,N5285,N5287,N5288,N5290,N5486 
	,N5532,N5538,N5539,N5542,N5543,N5546,N5553,N5556 
	,N5557,N5561,N5564,N5567,N5568,N5575,N5576,N5579 
	,N5580,N5583,N5587,N5588,N5591,N5594,N5595,N5596 
	,N5600,N5707,N5708,N5716,N5724,N5729,N5736,N5738 
	,N5743,N5746,N5754,N5857,N5869,N5875,N5893,N5912 
	,N5918,N5923,N5926,N5930,N5934,N5939,N5942,N5943 
	,N5947,N5953,N5956,N5961,N5966,N5969,N5973,N5978 
	,N5982,N5986,N5990,N5995,N5997,N5999,N6003,N6008 
	,N6011,N8056,N8072,N8080,N8086,N8092,N8098,N8139 
	,N8174,N8177,N8178,N8179,N8180,N8182,N8183,N8184 
	,N8185,N8186,N8188,N8194,N8202,N8208,N8222,N8229 
	,N8236,N8243,N8250,N8257,N13058,N13145,N13146,N13147 
	,N13148,N13149,N13150,N13151,N13152,N13268,N13269,N13272 
	,N13275,N13280,N13284,N13294,N13298,N13305,N13309,N13312 
	,N13314,N13350,N13352,N13354,N13359,N13362,N13365,N13366 
	,N13367,N13369,N13371,N13372,N13375,N13376,N13378,N13380 
	,N13384,N13385,N13387,N13388,N13389,N13392,N13433,N13439 
	,N13446,N13468,N13469,N13472,N13475,N13478,N13479,N13483 
	,N13485,N13486,N13489,N13493,N13499,N13500,N13503,N13504 
	,N13512,N13513,N13515,N13518,N13519,N13523,N13528,N13533 
	,N13535,N13540,N13593,N13596,N13597,N13599,N13601,N13604 
	,N13606,N13607,N13608,N13610,N13611,N13613,N13615,N13617 
	,N13621,N13627,N13629,N13634,N13635,N13681,N13683,N13685 
	,N13686,N13692,N13695,N13697,N13699,N13701,N13706,N13707 
	,N13710,N13719,N13722,N13730,N13732,N13734,N13738,N13740 
	,N13742,N13744,N13746,N13754,N13806,N13813,N13816,N13828 
	,N13835,N13842,N13849,N13856,N13858,N13864,N13872,N13877 
	,N13881,N13889,N13894,N13899,N13904,N13908,N13916;
XOR2XL cynw_cm_float_add2_ieee_I462 (.Y(inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
NAND2XL inst_cellmath__9_0_I463 (.Y(N3083), .A(a_exp[0]), .B(a_exp[1]));
AND4XL inst_cellmath__9_0_I8111 (.Y(N3085), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3138 (.Y(N8194), .A(a_exp[7]), .B(a_exp[6]), .C(N3085));
NOR2XL hyperpropagate_4_1_A_I3139 (.Y(inst_cellmath__9), .A(N3083), .B(N8194));
NOR2XL inst_cellmath__10__1__I476 (.Y(N3106), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__10__1__I477 (.Y(N3114), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__10__1__I478 (.Y(N3125), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__10__1__I479 (.Y(N3134), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__10__1__I8112 (.Y(N3119), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__10__1__I8113 (.Y(N3128), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__10__1__I8114 (.Y(N3138), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__10__1__I483 (.Y(N3123), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N3119));
NAND4XL inst_cellmath__10__1__I485 (.Y(N3117), .A(N3106), .B(N3125), .C(N3114), .D(N3134));
NOR4BX1 inst_cellmath__10__1__I8115 (.Y(inst_cellmath__10), .AN(N3123), .B(N3117), .C(N3128), .D(N3138));
NAND2XL inst_cellmath__14_0_I489 (.Y(N3168), .A(b_exp[0]), .B(b_exp[1]));
AND4XL inst_cellmath__14_0_I8116 (.Y(N3170), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3140 (.Y(N8202), .A(b_exp[7]), .B(b_exp[6]), .C(N3170));
NOR2XL hyperpropagate_4_1_A_I3141 (.Y(inst_cellmath__14), .A(N3168), .B(N8202));
NOR2XL inst_cellmath__15__3__I502 (.Y(N3191), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__15__3__I503 (.Y(N3199), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__15__3__I504 (.Y(N3210), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__15__3__I505 (.Y(N3219), .A(b_man[4]), .B(b_man[3]));
OR4X1 inst_cellmath__15__3__I8117 (.Y(N3204), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__15__3__I8118 (.Y(N3213), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__15__3__I8119 (.Y(N3223), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4X1 inst_cellmath__15__3__I509 (.Y(N3208), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N3204));
NAND4XL inst_cellmath__15__3__I511 (.Y(N3202), .A(N3191), .B(N3210), .C(N3199), .D(N3219));
NOR4BX1 inst_cellmath__15__3__I8120 (.Y(inst_cellmath__15), .AN(N3208), .B(N3202), .C(N3213), .D(N3223));
AND2XL inst_cellmath__59_0_I8068 (.Y(inst_cellmath__17), .A(inst_cellmath__14), .B(inst_cellmath__15));
AND2XL inst_cellmath__59_0_I8067 (.Y(inst_cellmath__12), .A(inst_cellmath__9), .B(inst_cellmath__10));
AND3XL cynw_cm_float_add2_ieee_I515 (.Y(N547), .A(inst_cellmath__17), .B(inst_cellmath__12), .C(inst_cellmath__39[25]));
NOR2BX1 cynw_cm_float_add2_ieee_I516 (.Y(inst_cellmath__13), .AN(inst_cellmath__9), .B(inst_cellmath__10));
NOR2BX1 cynw_cm_float_add2_ieee_I517 (.Y(inst_cellmath__18), .AN(inst_cellmath__14), .B(inst_cellmath__15));
OR4X1 inst_cellmath__11__2__I8121 (.Y(N3269), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 inst_cellmath__11__2__I8122 (.Y(N3273), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL inst_cellmath__11__2__I525 (.Y(inst_cellmath__11), .A(N3269), .B(N3273));
OR4X1 inst_cellmath__16__4__I8123 (.Y(N3291), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 inst_cellmath__16__4__I8124 (.Y(N3295), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL inst_cellmath__16__4__I532 (.Y(inst_cellmath__16), .A(N3291), .B(N3295));
NOR3BXL cynw_cm_float_add2_ieee_I534 (.Y(inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
CLKINVX8 cynw_cm_float_add2_ieee_I15 (.Y(N556), .A(b_exp[0]));
INVX2 cynw_cm_float_add2_ieee_I16 (.Y(N557), .A(b_exp[1]));
INVXL cynw_cm_float_add2_ieee_I17 (.Y(N558), .A(b_exp[2]));
INVXL cynw_cm_float_add2_ieee_I18 (.Y(N559), .A(b_exp[3]));
INVXL cynw_cm_float_add2_ieee_I19 (.Y(N560), .A(b_exp[4]));
INVXL cynw_cm_float_add2_ieee_I20 (.Y(N561), .A(b_exp[5]));
ADDHX1 inst_cellmath__28__8__I535 (.CO(N3321), .S(N565), .A(a_exp[0]), .B(N556));
ADDFHXL inst_cellmath__28__8__I536 (.CO(N3364), .S(N566), .A(N557), .B(a_exp[1]), .CI(N3321));
ADDFHXL inst_cellmath__28__8__I537 (.CO(N3338), .S(N567), .A(N558), .B(a_exp[2]), .CI(N3364));
ADDFHXL inst_cellmath__28__8__I538 (.CO(N3358), .S(N568), .A(N559), .B(a_exp[3]), .CI(N3338));
ADDFHXL inst_cellmath__28__8__I539 (.CO(N3331), .S(N569), .A(N560), .B(a_exp[4]), .CI(N3358));
ADDFHXL inst_cellmath__28__8__I540 (.CO(N3352), .S(N570), .A(N561), .B(a_exp[5]), .CI(N3331));
INVXL inst_cellmath__28__8__I8105 (.Y(N562), .A(b_exp[6]));
ADDFHXL inst_cellmath__28__8__I541 (.CO(N3324), .S(N571), .A(N562), .B(a_exp[6]), .CI(N3352));
NOR2X2 inst_cellmath__28__8__I2622 (.Y(N8056), .A(a_exp[0]), .B(N556));
INVX2 inst_cellmath__28__8__I2623 (.Y(N3333), .A(N8056));
ADDFHXL inst_cellmath__28__8__I546 (.CO(N3327), .S(inst_cellmath__27[1]), .A(N557), .B(a_exp[1]), .CI(N3333));
ADDFXL inst_cellmath__28__8__I547 (.CO(N3348), .S(inst_cellmath__27[2]), .A(N558), .B(a_exp[2]), .CI(N3327));
ADDFXL inst_cellmath__28__8__I548 (.CO(N3319), .S(inst_cellmath__27[3]), .A(N559), .B(a_exp[3]), .CI(N3348));
ADDFXL inst_cellmath__28__8__I549 (.CO(N3343), .S(inst_cellmath__27[4]), .A(N560), .B(a_exp[4]), .CI(N3319));
INVXL inst_cellmath__28__8__I8106 (.Y(N563), .A(b_exp[7]));
ADDFXL inst_cellmath__28__8__I8107 (.CO(N13816), .S(inst_cellmath__27[5]), .A(N561), .B(a_exp[5]), .CI(N3343));
ADDFXL inst_cellmath__28__8__I8108 (.CO(N13806), .S(inst_cellmath__27[6]), .A(N562), .B(a_exp[6]), .CI(N13816));
ADDFX1 inst_cellmath__28__8__I8109 (.CO(N13813), .S(inst_cellmath__27[7]), .A(N563), .B(a_exp[7]), .CI(N13806));
CLKINVX4 inst_cellmath__28__8__I8110 (.Y(inst_cellmath__27[8]), .A(N13813));
INVXL inst_cellmath__34_0_I554 (.Y(N3434), .A(a_man[1]));
INVXL inst_cellmath__34_0_I555 (.Y(N3501), .A(a_man[2]));
INVXL inst_cellmath__34_0_I556 (.Y(N3415), .A(a_man[3]));
INVXL inst_cellmath__34_0_I557 (.Y(N3480), .A(a_man[4]));
INVXL inst_cellmath__34_0_I558 (.Y(N3547), .A(a_man[5]));
INVXL inst_cellmath__34_0_I559 (.Y(N3461), .A(a_man[6]));
INVXL inst_cellmath__34_0_I560 (.Y(N3525), .A(a_man[7]));
INVXL inst_cellmath__34_0_I561 (.Y(N3444), .A(a_man[8]));
INVXL inst_cellmath__34_0_I562 (.Y(N3507), .A(a_man[9]));
INVXL inst_cellmath__34_0_I563 (.Y(N3421), .A(a_man[10]));
INVXL inst_cellmath__34_0_I564 (.Y(N3489), .A(a_man[11]));
INVXL inst_cellmath__34_0_I565 (.Y(N3405), .A(a_man[12]));
INVXL inst_cellmath__34_0_I566 (.Y(N3468), .A(a_man[13]));
INVXL inst_cellmath__34_0_I567 (.Y(N3535), .A(a_man[14]));
INVXL inst_cellmath__34_0_I568 (.Y(N3453), .A(a_man[15]));
INVXL inst_cellmath__34_0_I569 (.Y(N3515), .A(a_man[16]));
INVXL inst_cellmath__34_0_I570 (.Y(N3431), .A(a_man[17]));
INVXL inst_cellmath__34_0_I571 (.Y(N3498), .A(a_man[18]));
INVXL inst_cellmath__34_0_I572 (.Y(N3410), .A(a_man[19]));
INVXL inst_cellmath__34_0_I573 (.Y(N3478), .A(a_man[20]));
INVXL inst_cellmath__34_0_I574 (.Y(N3544), .A(a_man[21]));
INVXL inst_cellmath__34_0_I575 (.Y(N3457), .A(a_man[22]));
INVXL inst_cellmath__34_0_I576 (.Y(N3441), .A(b_man[0]));
NAND2XL inst_cellmath__34_0_I577 (.Y(N3449), .A(b_man[1]), .B(N3434));
NOR2XL inst_cellmath__34_0_I578 (.Y(N3414), .A(b_man[1]), .B(N3434));
NAND2XL inst_cellmath__34_0_I579 (.Y(N3546), .A(b_man[2]), .B(N3501));
NOR2XL inst_cellmath__34_0_I580 (.Y(N3512), .A(b_man[2]), .B(N3501));
NAND2XL inst_cellmath__34_0_I581 (.Y(N3494), .A(b_man[3]), .B(N3415));
NOR2XL inst_cellmath__34_0_I582 (.Y(N3460), .A(b_man[3]), .B(N3415));
NAND2XL inst_cellmath__34_0_I583 (.Y(N3443), .A(b_man[4]), .B(N3480));
NOR2XL inst_cellmath__34_0_I584 (.Y(N3408), .A(b_man[4]), .B(N3480));
NAND2XL inst_cellmath__34_0_I585 (.Y(N3540), .A(b_man[5]), .B(N3547));
NOR2XL inst_cellmath__34_0_I586 (.Y(N3506), .A(b_man[5]), .B(N3547));
NAND2XL inst_cellmath__34_0_I587 (.Y(N3488), .A(b_man[6]), .B(N3461));
NOR2XL inst_cellmath__34_0_I588 (.Y(N3455), .A(b_man[6]), .B(N3461));
NAND2XL inst_cellmath__34_0_I589 (.Y(N3437), .A(b_man[7]), .B(N3525));
NOR2XL inst_cellmath__34_0_I590 (.Y(N3404), .A(b_man[7]), .B(N3525));
NAND2XL inst_cellmath__34_0_I591 (.Y(N3534), .A(b_man[8]), .B(N3444));
NOR2XL inst_cellmath__34_0_I592 (.Y(N3503), .A(b_man[8]), .B(N3444));
NAND2XL inst_cellmath__34_0_I593 (.Y(N3483), .A(b_man[9]), .B(N3507));
NOR2XL inst_cellmath__34_0_I594 (.Y(N3451), .A(b_man[9]), .B(N3507));
NAND2XL inst_cellmath__34_0_I595 (.Y(N3430), .A(b_man[10]), .B(N3421));
NOR2XL inst_cellmath__34_0_I596 (.Y(N3550), .A(b_man[10]), .B(N3421));
NAND2XL inst_cellmath__34_0_I597 (.Y(N3528), .A(b_man[11]), .B(N3489));
NOR2XL inst_cellmath__34_0_I598 (.Y(N3496), .A(b_man[11]), .B(N3489));
NAND2XL inst_cellmath__34_0_I599 (.Y(N3477), .A(b_man[12]), .B(N3405));
NOR2XL inst_cellmath__34_0_I600 (.Y(N3446), .A(b_man[12]), .B(N3405));
NAND2XL inst_cellmath__34_0_I601 (.Y(N3424), .A(b_man[13]), .B(N3468));
NOR2XL inst_cellmath__34_0_I602 (.Y(N3542), .A(b_man[13]), .B(N3468));
NAND2XL inst_cellmath__34_0_I603 (.Y(N3524), .A(b_man[14]), .B(N3535));
NOR2XL inst_cellmath__34_0_I604 (.Y(N3492), .A(b_man[14]), .B(N3535));
NAND2XL inst_cellmath__34_0_I605 (.Y(N3471), .A(b_man[15]), .B(N3453));
NOR2XL inst_cellmath__34_0_I606 (.Y(N3439), .A(b_man[15]), .B(N3453));
NAND2XL inst_cellmath__34_0_I607 (.Y(N3419), .A(b_man[16]), .B(N3515));
NOR2XL inst_cellmath__34_0_I608 (.Y(N3537), .A(b_man[16]), .B(N3515));
NAND2XL inst_cellmath__34_0_I609 (.Y(N3518), .A(b_man[17]), .B(N3431));
NOR2XL inst_cellmath__34_0_I610 (.Y(N3485), .A(b_man[17]), .B(N3431));
NAND2XL inst_cellmath__34_0_I611 (.Y(N3465), .A(b_man[18]), .B(N3498));
NOR2XL inst_cellmath__34_0_I612 (.Y(N3433), .A(b_man[18]), .B(N3498));
NAND2XL inst_cellmath__34_0_I613 (.Y(N3413), .A(b_man[19]), .B(N3410));
NOR2XL inst_cellmath__34_0_I614 (.Y(N3530), .A(b_man[19]), .B(N3410));
NAND2XL inst_cellmath__34_0_I615 (.Y(N3511), .A(b_man[20]), .B(N3478));
NOR2XL inst_cellmath__34_0_I616 (.Y(N3479), .A(b_man[20]), .B(N3478));
NAND2XL inst_cellmath__34_0_I617 (.Y(N3459), .A(b_man[21]), .B(N3544));
NOR2XL inst_cellmath__34_0_I618 (.Y(N3426), .A(b_man[21]), .B(N3544));
OR2XL inst_cellmath__34_0_I619 (.Y(N3475), .A(b_man[22]), .B(N3457));
OAI21XL inst_cellmath__34_0_I620 (.Y(N3473), .A0(N3426), .A1(N3511), .B0(N3459));
NOR2XL inst_cellmath__34_0_I621 (.Y(N3505), .A(N3426), .B(N3479));
OAI21XL inst_cellmath__34_0_I622 (.Y(N3539), .A0(N3530), .A1(N3465), .B0(N3413));
NOR2XL inst_cellmath__34_0_I623 (.Y(N3420), .A(N3530), .B(N3433));
OAI21XL inst_cellmath__34_0_I624 (.Y(N3454), .A0(N3485), .A1(N3419), .B0(N3518));
NOR2XL inst_cellmath__34_0_I625 (.Y(N3487), .A(N3485), .B(N3537));
OAI21XL inst_cellmath__34_0_I626 (.Y(N3520), .A0(N3439), .A1(N3524), .B0(N3471));
NOR2XL inst_cellmath__34_0_I627 (.Y(N3403), .A(N3439), .B(N3492));
OAI21XL inst_cellmath__34_0_I628 (.Y(N3436), .A0(N3542), .A1(N3477), .B0(N3424));
NOR2XL inst_cellmath__34_0_I629 (.Y(N3467), .A(N3542), .B(N3446));
OAI21XL inst_cellmath__34_0_I630 (.Y(N3502), .A0(N3496), .A1(N3430), .B0(N3528));
NOR2XL inst_cellmath__34_0_I631 (.Y(N3532), .A(N3496), .B(N3550));
OAI21XL inst_cellmath__34_0_I632 (.Y(N3416), .A0(N3451), .A1(N3534), .B0(N3483));
OAI21XL inst_cellmath__34_0_I634 (.Y(N3482), .A0(N3404), .A1(N3488), .B0(N3437));
NOR2XL inst_cellmath__34_0_I635 (.Y(N3513), .A(N3404), .B(N3455));
OAI21XL inst_cellmath__34_0_I636 (.Y(N3548), .A0(N3506), .A1(N3443), .B0(N3540));
NOR2XL inst_cellmath__34_0_I637 (.Y(N3428), .A(N3506), .B(N3408));
OAI21XL inst_cellmath__34_0_I638 (.Y(N3462), .A0(N3460), .A1(N3546), .B0(N3494));
NOR2XL inst_cellmath__34_0_I639 (.Y(N3495), .A(N3460), .B(N3512));
OAI31X1 inst_cellmath__34_0_I640 (.Y(N3527), .A0(N3441), .A1(a_man[0]), .A2(N3414), .B0(N3449));
AOI22XL inst_cellmath__34_0_I641 (.Y(N3508), .A0(N3475), .A1(N3473), .B0(b_man[22]), .B1(N3457));
NAND2XL inst_cellmath__34_0_I642 (.Y(N3541), .A(N3475), .B(N3505));
AOI21XL inst_cellmath__34_0_I643 (.Y(N3423), .A0(N3420), .A1(N3454), .B0(N3539));
AOI21XL inst_cellmath__34_0_I644 (.Y(N3490), .A0(N3403), .A1(N3436), .B0(N3520));
NAND2XL inst_cellmath__34_0_I645 (.Y(N3522), .A(N3403), .B(N3467));
AOI21XL inst_cellmath__34_0_I646 (.Y(N3406), .A0(N3532), .A1(N3416), .B0(N3502));
NOR4BX1 inst_cellmath__34_0_I8126 (.Y(N3551), .AN(N3532), .B(N3451), .C(N3522), .D(N3503));
AOI21XL inst_cellmath__34_0_I648 (.Y(N3470), .A0(N3513), .A1(N3548), .B0(N3482));
NAND2XL inst_cellmath__34_0_I649 (.Y(N3504), .A(N3513), .B(N3428));
AOI21XL inst_cellmath__34_0_I650 (.Y(N3536), .A0(N3495), .A1(N3527), .B0(N3462));
NAND3BXL inst_cellmath__34_0_I651 (.Y(N3447), .AN(N3541), .B(N3420), .C(N3487));
OAI21XL inst_cellmath__34_0_I652 (.Y(N3517), .A0(N3522), .A1(N3406), .B0(N3490));
OAI21XL inst_cellmath__34_0_I654 (.Y(N3432), .A0(N3504), .A1(N3536), .B0(N3470));
AOI21XL inst_cellmath__34_0_I655 (.Y(N3499), .A0(N3551), .A1(N3432), .B0(N3517));
OA21X1 inst_cellmath__34_0_I656 (.Y(N3412), .A0(N3541), .A1(N3423), .B0(N3508));
OAI21XL inst_cellmath__34_0_I657 (.Y(inst_cellmath__34), .A0(N3447), .A1(N3499), .B0(N3412));
ADDFHXL inst_cellmath__59_0_I7917 (.CO(N3367), .S(N572), .A(N563), .B(a_exp[7]), .CI(N3324));
NOR2BX2 cynw_cm_float_add2_ieee_I658 (.Y(N575), .AN(inst_cellmath__34), .B(N3367));
NOR2X6 cynw_cm_float_add2_ieee_I659 (.Y(inst_cellmath__32), .A(inst_cellmath__27[8]), .B(N575));
MX2XL cynw_cm_float_add2_ieee_I660 (.Y(inst_cellmath__48), .A(b_sign), .B(a_sign), .S0(inst_cellmath__32));
XOR2XL inst_cellmath__35_0_I2967 (.Y(N3682), .A(N556), .B(a_exp[0]));
INVXL inst_cellmath__35_0_I662 (.Y(N3691), .A(inst_cellmath__27[1]));
INVXL inst_cellmath__35_0_I663 (.Y(N3698), .A(inst_cellmath__27[2]));
INVXL inst_cellmath__35_0_I664 (.Y(N3671), .A(inst_cellmath__27[3]));
INVXL inst_cellmath__35_0_I665 (.Y(N3678), .A(inst_cellmath__27[4]));
INVXL inst_cellmath__35_0_I666 (.Y(N3686), .A(inst_cellmath__27[5]));
INVXL inst_cellmath__35_0_I667 (.Y(N3694), .A(inst_cellmath__27[6]));
INVXL inst_cellmath__35_0_I668 (.Y(N3701), .A(inst_cellmath__27[7]));
INVX3 inst_cellmath__35_0_I669 (.Y(N3688), .A(inst_cellmath__27[8]));
AOI22X2 inst_cellmath__35_0_I670 (.Y(inst_cellmath__35[0]), .A0(N3682), .A1(N3688), .B0(N565), .B1(inst_cellmath__27[8]));
AOI22X1 inst_cellmath__35_0_I671 (.Y(inst_cellmath__35[1]), .A0(N3691), .A1(N3688), .B0(N566), .B1(inst_cellmath__27[8]));
AOI22X2 inst_cellmath__35_0_I672 (.Y(inst_cellmath__35[2]), .A0(N3698), .A1(N3688), .B0(N567), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I673 (.Y(inst_cellmath__35[3]), .A0(N3671), .A1(N3688), .B0(N568), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I674 (.Y(inst_cellmath__35[4]), .A0(N3678), .A1(N3688), .B0(N569), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I675 (.Y(inst_cellmath__35[5]), .A0(N3686), .A1(N3688), .B0(N570), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I676 (.Y(inst_cellmath__35[6]), .A0(N3694), .A1(N3688), .B0(N571), .B1(inst_cellmath__27[8]));
AOI22XL inst_cellmath__35_0_I677 (.Y(inst_cellmath__35[7]), .A0(N3688), .A1(N3701), .B0(N572), .B1(inst_cellmath__27[8]));
OAI211X1 inst_cellmath__30_0_I678 (.Y(N3730), .A0(inst_cellmath__35[1]), .A1(inst_cellmath__35[2]), .B0(inst_cellmath__35[4]), .C0(inst_cellmath__35[3]));
NOR3BX1 inst_cellmath__30_0_I679 (.Y(N3729), .AN(N3730), .B(inst_cellmath__35[6]), .C(inst_cellmath__35[5]));
NAND2BX2 inst_cellmath__30_0_I680 (.Y(inst_cellmath__30), .AN(inst_cellmath__35[7]), .B(N3729));
OR2X1 cynw_cm_float_add2_ieee_I681 (.Y(inst_cellmath__31), .A(inst_cellmath__11), .B(inst_cellmath__16));
INVX12 inst_cellmath__36__15__I684 (.Y(N3769), .A(inst_cellmath__32));
INVX1 inst_cellmath__36__15__I7655 (.Y(N13145), .A(N3769));
INVXL inst_cellmath__36__15__I7885 (.Y(N13150), .A(N13145));
MX2XL inst_cellmath__36__15__I7886 (.Y(N13366), .A(a_man[1]), .B(b_man[1]), .S0(N13150));
MXI2XL inst_cellmath__36__15__I7887 (.Y(N13384), .A(a_man[2]), .B(b_man[2]), .S0(N13150));
MX2XL inst_cellmath__36__15__I7888 (.Y(N13376), .A(a_man[2]), .B(b_man[2]), .S0(N13150));
NOR2X2 inst_cellmath__33_49_24_I2973 (.Y(N4277), .A(inst_cellmath__31), .B(inst_cellmath__30));
INVX3 inst_cellmath__37_0_I846 (.Y(N3842), .A(inst_cellmath__35[3]));
CLKINVX8 inst_cellmath__37_0_I847 (.Y(N3890), .A(N3842));
INVX2 inst_cellmath__37_0_I797 (.Y(N3920), .A(inst_cellmath__35[4]));
CLKINVX6 inst_cellmath__37_0_I798 (.Y(N3964), .A(N3920));
CLKINVX12 inst_cellmath__37_0_I764 (.Y(N3992), .A(inst_cellmath__35[1]));
CLKINVX4 inst_cellmath__37_0_I765 (.Y(N4041), .A(N3992));
INVX4 inst_cellmath__37_0_I708 (.Y(N4021), .A(inst_cellmath__35[0]));
CLKINVX6 inst_cellmath__37_0_I733 (.Y(N3851), .A(inst_cellmath__35[2]));
NAND2XL inst_cellmath__37_0_I763 (.Y(N3960), .A(N4021), .B(N3851));
NOR2XL inst_cellmath__37_0_I796 (.Y(N4037), .A(N3960), .B(N4041));
CLKINVX8 inst_cellmath__37_0_I734 (.Y(N3901), .A(N3851));
MX2XL inst_cellmath__36__15__I697 (.Y(inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(N3769));
MXI2XL mx2a_A_I8269 (.Y(N13828), .A(b_man[11]), .B(a_man[11]), .S0(N3769));
INVXL mx2a_A_I8270 (.Y(inst_cellmath__36[37]), .A(N13828));
MX2XL inst_cellmath__37_0_I721 (.Y(N3858), .A(inst_cellmath__36[38]), .B(inst_cellmath__36[37]), .S0(N4021));
MX2XL inst_cellmath__36__15__I693 (.Y(inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(N3769));
MX2XL inst_cellmath__36__15__I692 (.Y(inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(N3769));
MX2XL inst_cellmath__37_0_I717 (.Y(N3884), .A(inst_cellmath__36[34]), .B(inst_cellmath__36[33]), .S0(N4021));
AOI22X1 inst_cellmath__37_0_I747 (.Y(N3932), .A0(N3858), .A1(N3901), .B0(N3884), .B1(N3851));
MXI2XL mx2a_A_I8271 (.Y(N13835), .A(b_man[14]), .B(a_man[14]), .S0(N3769));
INVXL mx2a_A_I8272 (.Y(inst_cellmath__36[40]), .A(N13835));
MXI2XL mx2a_A_I8273 (.Y(N13842), .A(b_man[13]), .B(a_man[13]), .S0(N3769));
INVXL mx2a_A_I8274 (.Y(inst_cellmath__36[39]), .A(N13842));
MX2XL inst_cellmath__37_0_I723 (.Y(N3950), .A(inst_cellmath__36[40]), .B(inst_cellmath__36[39]), .S0(N4021));
MX2XL inst_cellmath__36__15__I2971 (.Y(inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(N3769));
MX2XL inst_cellmath__36__15__I2970 (.Y(inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(N3769));
MX2XL inst_cellmath__37_0_I719 (.Y(N3979), .A(inst_cellmath__36[36]), .B(inst_cellmath__36[35]), .S0(N4021));
AOI22X1 inst_cellmath__37_0_I749 (.Y(N4024), .A0(N3901), .A1(N3950), .B0(N3979), .B1(N3851));
AOI22XL inst_cellmath__37_0_I780 (.Y(N4055), .A0(N3992), .A1(N3932), .B0(N4041), .B1(N4024));
AOI22XL inst_cellmath__37_0_I829 (.Y(N4042), .A0(N4037), .A1(N3964), .B0(N3920), .B1(N4055));
MX2XL inst_cellmath__36__15__I685 (.Y(inst_cellmath__36[26]), .A(b_man[0]), .B(a_man[0]), .S0(N3769));
NOR2BX1 inst_cellmath__37_0_I709 (.Y(N3892), .AN(inst_cellmath__36[26]), .B(N4021));
MXI2XL mx2a_A_I7575 (.Y(N13058), .A(b_man[4]), .B(a_man[4]), .S0(N3769));
INVXL mx2a_A_I7576 (.Y(inst_cellmath__36[30]), .A(N13058));
MXI2XL mx2a_A_I8275 (.Y(N13849), .A(b_man[3]), .B(a_man[3]), .S0(N3769));
INVXL mx2a_A_I8276 (.Y(inst_cellmath__36[29]), .A(N13849));
MX2XL inst_cellmath__37_0_I713 (.Y(N3915), .A(inst_cellmath__36[30]), .B(inst_cellmath__36[29]), .S0(N4021));
AOI22X1 inst_cellmath__37_0_I2760 (.Y(N3983), .A0(N3851), .A1(N3892), .B0(N3901), .B1(N3915));
MX2XL inst_cellmath__36__15__I2969 (.Y(inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(N3769));
MX2XL inst_cellmath__36__15__I8129 (.Y(inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(N3769));
MX2X1 inst_cellmath__37_0_I715 (.Y(N4006), .A(inst_cellmath__36[32]), .B(inst_cellmath__36[31]), .S0(N4021));
MX2XL inst_cellmath__36__15__I687 (.Y(inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(N3769));
MX2XL inst_cellmath__36__15__I686 (.Y(inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(N3769));
MX2X1 inst_cellmath__37_0_I711 (.Y(N4033), .A(inst_cellmath__36[28]), .B(inst_cellmath__36[27]), .S0(N4021));
AOI22X2 inst_cellmath__37_0_I741 (.Y(N3864), .A0(N3901), .A1(N4006), .B0(N4033), .B1(N3851));
AOI22X1 inst_cellmath__37_0_I772 (.Y(N3891), .A0(N3992), .A1(N3983), .B0(N4041), .B1(N3864));
MX2XL inst_cellmath__36__15__I705 (.Y(inst_cellmath__36[46]), .A(b_man[20]), .B(a_man[20]), .S0(N3769));
MX2XL inst_cellmath__36__15__I704 (.Y(inst_cellmath__36[45]), .A(b_man[19]), .B(a_man[19]), .S0(N3769));
MX2XL inst_cellmath__37_0_I729 (.Y(N4017), .A(inst_cellmath__36[46]), .B(inst_cellmath__36[45]), .S0(N4021));
MX2XL inst_cellmath__36__15__I701 (.Y(inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(N3769));
MX2XL inst_cellmath__36__15__I700 (.Y(inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(N3769));
MX2XL inst_cellmath__37_0_I725 (.Y(N4047), .A(inst_cellmath__36[42]), .B(inst_cellmath__36[41]), .S0(N4021));
AOI22XL inst_cellmath__37_0_I755 (.Y(N3874), .A0(N3901), .A1(N4017), .B0(N4047), .B1(N3851));
MX2XL inst_cellmath__36__15__I707 (.Y(inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(N3769));
MX2XL inst_cellmath__36__15__I706 (.Y(inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(N3769));
MX2XL inst_cellmath__37_0_I731 (.Y(N3896), .A(inst_cellmath__36[48]), .B(inst_cellmath__36[47]), .S0(N4021));
MX2XL inst_cellmath__36__15__I703 (.Y(inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(N3769));
MX2XL inst_cellmath__36__15__I702 (.Y(inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(N3769));
MX2XL inst_cellmath__37_0_I727 (.Y(N3926), .A(inst_cellmath__36[44]), .B(inst_cellmath__36[43]), .S0(N4021));
AOI22X1 inst_cellmath__37_0_I757 (.Y(N3968), .A0(N3901), .A1(N3896), .B0(N3926), .B1(N3851));
AOI22XL inst_cellmath__37_0_I788 (.Y(N3998), .A0(N3992), .A1(N3874), .B0(N4041), .B1(N3968));
AOI22X1 inst_cellmath__37_0_I2764 (.Y(N3879), .A0(N3891), .A1(N3920), .B0(N3964), .B1(N3998));
AOI22XL inst_cellmath__37_0_I2714 (.Y(inst_cellmath__37[25]), .A0(N3890), .A1(N4042), .B0(N3842), .B1(N3879));
AND2XL inst_cellmath__33_49_24_I900 (.Y(inst_cellmath__33[25]), .A(N4277), .B(inst_cellmath__37[25]));
INVX1 inst_cellmath__36__15__I8036 (.Y(N4400), .A(inst_cellmath__39[25]));
XNOR2X1 inst_cellmath__39__19__2mx_I973 (.Y(inst_cellmath__39[0]), .A(N4400), .B(inst_cellmath__33[25]));
MX2XL inst_cellmath__37_0_I728 (.Y(N3971), .A(inst_cellmath__36[45]), .B(inst_cellmath__36[44]), .S0(N4021));
MX2XL inst_cellmath__37_0_I724 (.Y(N3999), .A(inst_cellmath__36[41]), .B(inst_cellmath__36[40]), .S0(N4021));
AOI22X1 inst_cellmath__37_0_I754 (.Y(N4044), .A0(N3901), .A1(N3971), .B0(N3851), .B1(N3999));
MX2XL inst_cellmath__37_0_I730 (.Y(N3849), .A(inst_cellmath__36[47]), .B(inst_cellmath__36[46]), .S0(N4021));
MX2X1 inst_cellmath__37_0_I726 (.Y(N3877), .A(inst_cellmath__36[43]), .B(inst_cellmath__36[42]), .S0(N4021));
AOI22X2 inst_cellmath__37_0_I756 (.Y(N3923), .A0(N3901), .A1(N3849), .B0(N3851), .B1(N3877));
AOI22X1 inst_cellmath__37_0_I787 (.Y(N3949), .A0(N3992), .A1(N4044), .B0(N4041), .B1(N3923));
MX2XL inst_cellmath__37_0_I712 (.Y(N3867), .A(inst_cellmath__36[29]), .B(inst_cellmath__36[28]), .S0(N4021));
NAND2XL inst_cellmath__37_0_I738 (.Y(N3889), .A(N3901), .B(N3867));
MX2XL inst_cellmath__37_0_I714 (.Y(N3959), .A(inst_cellmath__36[31]), .B(inst_cellmath__36[30]), .S0(N4021));
MX2XL inst_cellmath__37_0_I710 (.Y(N3985), .A(inst_cellmath__36[27]), .B(inst_cellmath__36[26]), .S0(N4021));
AOI22X2 inst_cellmath__37_0_I740 (.Y(N4031), .A0(N3901), .A1(N3959), .B0(N3985), .B1(N3851));
AOI22XL inst_cellmath__37_0_I771 (.Y(N3843), .A0(N3889), .A1(N3992), .B0(N4041), .B1(N4031));
AOI22XL inst_cellmath__37_0_I820 (.Y(N4051), .A0(N3964), .A1(N3949), .B0(N3843), .B1(N3920));
NAND2BXL inst_cellmath__37_0_I732 (.Y(N3942), .AN(inst_cellmath__36[48]), .B(N4021));
NAND2XL inst_cellmath__37_0_I762 (.Y(N3868), .A(N3942), .B(N3851));
NOR2XL inst_cellmath__37_0_I795 (.Y(N3895), .A(N3868), .B(N4041));
MX2XL inst_cellmath__37_0_I720 (.Y(N4027), .A(inst_cellmath__36[37]), .B(inst_cellmath__36[36]), .S0(N4021));
MX2XL inst_cellmath__37_0_I716 (.Y(N4056), .A(inst_cellmath__36[33]), .B(inst_cellmath__36[32]), .S0(N4021));
AOI22X1 inst_cellmath__37_0_I746 (.Y(N3881), .A0(N3901), .A1(N4027), .B0(N3851), .B1(N4056));
MX2XL inst_cellmath__37_0_I722 (.Y(N3907), .A(inst_cellmath__36[39]), .B(inst_cellmath__36[38]), .S0(N4021));
MX2XL inst_cellmath__37_0_I718 (.Y(N3935), .A(inst_cellmath__36[35]), .B(inst_cellmath__36[34]), .S0(N4021));
AOI22X1 inst_cellmath__37_0_I748 (.Y(N3975), .A0(N3907), .A1(N3901), .B0(N3851), .B1(N3935));
AOI22XL inst_cellmath__37_0_I779 (.Y(N4005), .A0(N3881), .A1(N3992), .B0(N4041), .B1(N3975));
AOI22XL inst_cellmath__37_0_I828 (.Y(N3994), .A0(N3895), .A1(N3964), .B0(N3920), .B1(N4005));
AOI22XL inst_cellmath__37_0_I872 (.Y(inst_cellmath__37[24]), .A0(N3842), .A1(N4051), .B0(N3994), .B1(N3890));
AND2XL inst_cellmath__33_49_24_I899 (.Y(inst_cellmath__33[24]), .A(inst_cellmath__37[24]), .B(N4277));
AOI22X1 inst_cellmath__37_0_I743 (.Y(N3956), .A0(N3884), .A1(N3901), .B0(N3851), .B1(N3915));
AOI22XL inst_cellmath__37_0_I774 (.Y(N3984), .A0(N3992), .A1(N3864), .B0(N4041), .B1(N3956));
NAND2XL inst_cellmath__37_0_I807 (.Y(N3928), .A(N3964), .B(N3984));
AOI22X1 inst_cellmath__37_0_I751 (.Y(N3904), .A0(N3901), .A1(N4047), .B0(N3858), .B1(N3851));
AOI22X2 inst_cellmath__37_0_I782 (.Y(N3934), .A0(N3992), .A1(N4024), .B0(N4041), .B1(N3904));
NAND2XL inst_cellmath__37_0_I735 (.Y(N4040), .A(N3901), .B(N3892));
NOR2XL inst_cellmath__37_0_I766 (.Y(N3852), .A(N3992), .B(N4040));
AOI22X2 inst_cellmath__37_0_I815 (.Y(N4029), .A0(N3964), .A1(N3934), .B0(N3852), .B1(N3920));
AOI22XL inst_cellmath__37_0_I859 (.Y(inst_cellmath__37[11]), .A0(N3842), .A1(N3928), .B0(N4029), .B1(N3890));
AOI22XL inst_cellmath__37_0_I745 (.Y(N4053), .A0(N3901), .A1(N3979), .B0(N4006), .B1(N3851));
AOI22XL inst_cellmath__37_0_I778 (.Y(N3958), .A0(N3992), .A1(N4053), .B0(N4041), .B1(N3932));
NAND2XL inst_cellmath__37_0_I811 (.Y(N3869), .A(N3964), .B(N3958));
NAND2XL inst_cellmath__37_0_I737 (.Y(N4011), .A(N3901), .B(N4033));
AOI22XL inst_cellmath__37_0_I770 (.Y(N4012), .A0(N4011), .A1(N3992), .B0(N4041), .B1(N3983));
AOI22XL inst_cellmath__37_0_I2655 (.Y(N3996), .A0(N3851), .A1(N3950), .B0(N3926), .B1(N3901));
AOI22XL inst_cellmath__37_0_I786 (.Y(N3906), .A0(N3992), .A1(N3996), .B0(N4041), .B1(N3874));
AOI22X1 inst_cellmath__37_0_I2763 (.Y(N4001), .A0(N4012), .A1(N3920), .B0(N3964), .B1(N3906));
AOI22XL inst_cellmath__37_0_I863 (.Y(inst_cellmath__37[15]), .A0(N3869), .A1(N3842), .B0(N3890), .B1(N4001));
AOI22XL inst_cellmath__37_0_I768 (.Y(N3921), .A0(N3992), .A1(N4040), .B0(N4041), .B1(N4011));
AOI22XL inst_cellmath__37_0_I2656 (.Y(N4026), .A0(N4041), .A1(N3996), .B0(N3992), .B1(N3904));
AOI22X1 inst_cellmath__37_0_I2658 (.Y(N3909), .A0(N3921), .A1(N3920), .B0(N3964), .B1(N4026));
AOI22XL inst_cellmath__37_0_I776 (.Y(N3866), .A0(N3992), .A1(N3956), .B0(N4041), .B1(N4053));
NAND2X1 inst_cellmath__37_0_I809 (.Y(N3899), .A(N3964), .B(N3866));
AOI22X1 inst_cellmath__37_0_I2660 (.Y(inst_cellmath__37[13]), .A0(N3890), .A1(N3909), .B0(N3842), .B1(N3899));
NAND2X1 inst_cellmath__37_0_I812 (.Y(N3962), .A(N3964), .B(N4005));
AOI22X1 inst_cellmath__37_0_I864 (.Y(inst_cellmath__37[16]), .A0(N3842), .A1(N3962), .B0(N3890), .B1(N4051));
NOR4X1 inst_cellmath__42__22__I937 (.Y(N4342), .A(inst_cellmath__37[11]), .B(inst_cellmath__37[16]), .C(inst_cellmath__37[15]), .D(inst_cellmath__37[13]));
AOI22X1 inst_cellmath__37_0_I750 (.Y(N3855), .A0(N3901), .A1(N3999), .B0(N3851), .B1(N4027));
AOI22XL inst_cellmath__37_0_I781 (.Y(N3883), .A0(N3992), .A1(N3975), .B0(N4041), .B1(N3855));
NAND2XL inst_cellmath__37_0_I814 (.Y(N3937), .A(N3964), .B(N3883));
AOI22XL inst_cellmath__37_0_I758 (.Y(N4014), .A0(N3942), .A1(N3901), .B0(N3851), .B1(N3971));
AOI22X1 inst_cellmath__37_0_I789 (.Y(N4046), .A0(N3992), .A1(N3923), .B0(N4041), .B1(N4014));
AOI22X1 inst_cellmath__37_0_I742 (.Y(N3911), .A0(N3901), .A1(N4056), .B0(N3851), .B1(N3867));
AOI22X1 inst_cellmath__37_0_I773 (.Y(N3939), .A0(N3992), .A1(N4031), .B0(N4041), .B1(N3911));
AOI22X1 inst_cellmath__37_0_I822 (.Y(N3930), .A0(N3964), .A1(N4046), .B0(N3920), .B1(N3939));
AOI22XL inst_cellmath__37_0_I866 (.Y(inst_cellmath__37[18]), .A0(N3937), .A1(N3842), .B0(N3890), .B1(N3930));
AOI22XL inst_cellmath__37_0_I744 (.Y(N4003), .A0(N3901), .A1(N3935), .B0(N3851), .B1(N3959));
AOI22XL inst_cellmath__37_0_I777 (.Y(N3913), .A0(N3992), .A1(N4003), .B0(N4041), .B1(N3881));
NAND2X1 inst_cellmath__37_0_I810 (.Y(N3990), .A(N3964), .B(N3913));
AOI22X2 inst_cellmath__37_0_I752 (.Y(N3947), .A0(N3901), .A1(N3877), .B0(N3851), .B1(N3907));
AOI22X1 inst_cellmath__37_0_I785 (.Y(N3857), .A0(N3992), .A1(N3947), .B0(N4041), .B1(N4044));
NAND2XL inst_cellmath__37_0_I736 (.Y(N3919), .A(N3901), .B(N3985));
AOI22XL inst_cellmath__37_0_I769 (.Y(N3965), .A0(N3919), .A1(N3992), .B0(N3889), .B1(N4041));
AOI22X1 inst_cellmath__37_0_I818 (.Y(N3954), .A0(N3964), .A1(N3857), .B0(N3920), .B1(N3965));
AOI22XL inst_cellmath__37_0_I862 (.Y(inst_cellmath__37[14]), .A0(N3990), .A1(N3842), .B0(N3890), .B1(N3954));
NAND2XL inst_cellmath__37_0_I799 (.Y(N4035), .A(N3964), .B(N3852));
AOI22X1 inst_cellmath__37_0_I851 (.Y(inst_cellmath__37[3]), .A0(N3842), .A1(N4035), .B0(N3890), .B1(N3928));
NAND2XL inst_cellmath__37_0_I803 (.Y(N3980), .A(N3964), .B(N4012));
AOI22XL inst_cellmath__37_0_I855 (.Y(inst_cellmath__37[7]), .A0(N3980), .A1(N3842), .B0(N3890), .B1(N3869));
NOR2X1 inst_cellmath__42__22__I928 (.Y(N4363), .A(inst_cellmath__37[3]), .B(inst_cellmath__37[7]));
NAND2XL inst_cellmath__37_0_I801 (.Y(N4008), .A(N3964), .B(N3921));
AOI22X1 inst_cellmath__37_0_I853 (.Y(inst_cellmath__37[5]), .A0(N4008), .A1(N3842), .B0(N3890), .B1(N3899));
NAND2X1 inst_cellmath__37_0_I805 (.Y(N3952), .A(N3964), .B(N3891));
NAND2X1 inst_cellmath__37_0_I813 (.Y(N3840), .A(N3964), .B(N4055));
AOI22XL inst_cellmath__37_0_I857 (.Y(inst_cellmath__37[9]), .A0(N3952), .A1(N3842), .B0(N3890), .B1(N3840));
NOR2X1 inst_cellmath__42__22__I929 (.Y(N4372), .A(inst_cellmath__37[5]), .B(inst_cellmath__37[9]));
NAND2X1 inst_cellmath__42__22__I934 (.Y(N4335), .A(N4363), .B(N4372));
NOR3X1 inst_cellmath__42__22__I938 (.Y(N4339), .A(inst_cellmath__37[18]), .B(inst_cellmath__37[14]), .C(N4335));
NAND2XL inst_cellmath__42__22__I941 (.Y(N4353), .A(N4339), .B(N4342));
NAND2XL inst_cellmath__37_0_I761 (.Y(N3986), .A(N3896), .B(N3851));
AOI22XL inst_cellmath__37_0_I794 (.Y(N3848), .A0(N3992), .A1(N3986), .B0(N3960), .B1(N4041));
AOI22XL inst_cellmath__37_0_I827 (.Y(N3945), .A0(N3848), .A1(N3964), .B0(N3920), .B1(N3958));
AOI22XL inst_cellmath__37_0_I871 (.Y(inst_cellmath__37[23]), .A0(N3842), .A1(N4001), .B0(N3945), .B1(N3890));
NAND2XL inst_cellmath__37_0_I760 (.Y(N3893), .A(N3851), .B(N3849));
AOI22XL inst_cellmath__37_0_I793 (.Y(N4016), .A0(N3893), .A1(N3992), .B0(N3868), .B1(N4041));
AOI22XL inst_cellmath__37_0_I826 (.Y(N3902), .A0(N4016), .A1(N3964), .B0(N3920), .B1(N3913));
AOI22X1 inst_cellmath__37_0_I870 (.Y(inst_cellmath__37[22]), .A0(N3842), .A1(N3954), .B0(N3890), .B1(N3902));
NAND2X1 inst_cellmath__37_0_I804 (.Y(N3860), .A(N3964), .B(N3843));
AOI22X1 inst_cellmath__37_0_I856 (.Y(inst_cellmath__37[8]), .A0(N3860), .A1(N3842), .B0(N3890), .B1(N3962));
NAND2XL inst_cellmath__37_0_I802 (.Y(N3886), .A(N3965), .B(N3964));
AOI22X1 inst_cellmath__37_0_I854 (.Y(inst_cellmath__37[6]), .A0(N3842), .A1(N3886), .B0(N3890), .B1(N3990));
NOR2X1 inst_cellmath__42__22__I930 (.Y(N4337), .A(inst_cellmath__37[8]), .B(inst_cellmath__37[6]));
NOR2XL inst_cellmath__37_0_I767 (.Y(N3993), .A(N3919), .B(N3992));
NAND2X1 inst_cellmath__37_0_I800 (.Y(N3916), .A(N3964), .B(N3993));
AOI22X1 inst_cellmath__37_0_I775 (.Y(N4032), .A0(N3992), .A1(N3911), .B0(N4041), .B1(N4003));
NAND2X1 inst_cellmath__37_0_I808 (.Y(N4019), .A(N3964), .B(N4032));
AOI22X1 inst_cellmath__37_0_I852 (.Y(inst_cellmath__37[4]), .A0(N3916), .A1(N3842), .B0(N4019), .B1(N3890));
NAND2X1 inst_cellmath__37_0_I806 (.Y(N4049), .A(N3964), .B(N3939));
AOI22XL inst_cellmath__37_0_I858 (.Y(inst_cellmath__37[10]), .A0(N3842), .A1(N4049), .B0(N3890), .B1(N3937));
NOR2X1 inst_cellmath__42__22__I931 (.Y(N4346), .A(inst_cellmath__37[4]), .B(inst_cellmath__37[10]));
NAND2X1 inst_cellmath__42__22__I935 (.Y(N4349), .A(N4337), .B(N4346));
NOR3X1 inst_cellmath__42__22__I939 (.Y(N4362), .A(inst_cellmath__37[23]), .B(inst_cellmath__37[22]), .C(N4349));
AOI22X2 inst_cellmath__37_0_I783 (.Y(N3977), .A0(N3992), .A1(N3855), .B0(N4041), .B1(N3947));
AOI22X2 inst_cellmath__37_0_I816 (.Y(N3862), .A0(N3964), .A1(N3977), .B0(N3993), .B1(N3920));
AOI22X1 inst_cellmath__37_0_I791 (.Y(N3925), .A0(N3992), .A1(N4014), .B0(N4041), .B1(N3893));
AOI22XL inst_cellmath__37_0_I824 (.Y(N4022), .A0(N3964), .A1(N3925), .B0(N3920), .B1(N4032));
AOI22XL inst_cellmath__37_0_I868 (.Y(inst_cellmath__37[20]), .A0(N3842), .A1(N3862), .B0(N4022), .B1(N3890));
AOI22XL inst_cellmath__37_0_I759 (.Y(N3846), .A0(N4021), .A1(N3901), .B0(N3851), .B1(N4017));
AOI22XL inst_cellmath__37_0_I792 (.Y(N3970), .A0(N3992), .A1(N3846), .B0(N3986), .B1(N4041));
AOI22XL inst_cellmath__37_0_I825 (.Y(N3853), .A0(N3964), .A1(N3970), .B0(N3920), .B1(N3866));
AOI22XL inst_cellmath__37_0_I2662 (.Y(inst_cellmath__37[21]), .A0(N3890), .A1(N3853), .B0(N3842), .B1(N3909));
AOI22X2 inst_cellmath__37_0_I860 (.Y(inst_cellmath__37[12]), .A0(N3842), .A1(N4019), .B0(N3890), .B1(N3862));
AOI22X1 inst_cellmath__37_0_I865 (.Y(inst_cellmath__37[17]), .A0(N3842), .A1(N3840), .B0(N3890), .B1(N3879));
NOR2X1 inst_cellmath__42__22__I932 (.Y(N4366), .A(inst_cellmath__37[12]), .B(inst_cellmath__37[17]));
NOR2X1 inst_cellmath__37_0_I848 (.Y(inst_cellmath__37[0]), .A(N3842), .B(N3860));
NOR2X1 inst_cellmath__42__22__I925 (.Y(N4333), .A(inst_cellmath__30), .B(inst_cellmath__37[0]));
INVXL gena_A_I8277 (.Y(N13856), .A(N3842));
NAND2XL gena_A_I8278 (.Y(N13858), .A(N3952), .B(N4049));
NAND2XL gena_A_I8279 (.Y(N4343), .A(N13856), .B(N13858));
NAND2X1 inst_cellmath__42__22__I927 (.Y(N4354), .A(N4333), .B(N4343));
AOI22X1 inst_cellmath__37_0_I2709 (.Y(N3876), .A0(N4041), .A1(N3846), .B0(N3992), .B1(N3968));
AOI22XL inst_cellmath__37_0_I823 (.Y(N3973), .A0(N3964), .A1(N3876), .B0(N3920), .B1(N3984));
AOI22X1 inst_cellmath__37_0_I867 (.Y(inst_cellmath__37[19]), .A0(N3842), .A1(N4029), .B0(N3890), .B1(N3973));
NOR2X1 inst_cellmath__42__22__I933 (.Y(N4351), .A(N4354), .B(inst_cellmath__37[19]));
NAND2X1 inst_cellmath__42__22__I936 (.Y(N4356), .A(N4366), .B(N4351));
NOR3X1 inst_cellmath__42__22__I940 (.Y(N4332), .A(inst_cellmath__37[20]), .B(inst_cellmath__37[21]), .C(N4356));
NAND2X1 inst_cellmath__42__22__I942 (.Y(N4371), .A(N4362), .B(N4332));
AOI2BB1X2 cynw_cm_float_add2_ieee_I7465 (.Y(inst_cellmath__42), .A0N(N4353), .A1N(N4371), .B0(inst_cellmath__31));
NOR3X2 cynw_cm_float_add2_ieee_I946 (.Y(inst_cellmath__44), .A(inst_cellmath__33[24]), .B(N4400), .C(inst_cellmath__42));
NAND2X2 inst_cellmath__36__15__I7889 (.Y(N13375), .A(inst_cellmath__39[0]), .B(inst_cellmath__44));
MXI2XL cynw_cm_float_add2_ieee_I949 (.Y(N655), .A(a_man[0]), .B(b_man[0]), .S0(N13150));
NAND2XL inst_cellmath__37_0_I830 (.Y(N3872), .A(N3920), .B(N3883));
AOI22X1 inst_cellmath__37_0_I874 (.Y(inst_cellmath__37[26]), .A0(N3842), .A1(N3930), .B0(N3872), .B1(N3890));
NAND2X1 inst_cellmath__33_49_24_I901 (.Y(inst_cellmath__33[26]), .A(N4277), .B(inst_cellmath__37[26]));
INVXL xnor2_A_I8280 (.Y(N13864), .A(N4400));
MXI2XL xnor2_A_I8281 (.Y(inst_cellmath__39[1]), .A(N4400), .B(N13864), .S0(inst_cellmath__33[26]));
NAND2XL inst_cellmath__36__15__I7890 (.Y(N13352), .A(N655), .B(inst_cellmath__39[1]));
XOR2X1 inst_cellmath__36__15__I7891 (.Y(N13388), .A(N655), .B(inst_cellmath__39[1]));
NAND2XL inst_cellmath__37_0_I831 (.Y(N3966), .A(N3934), .B(N3920));
AOI22XL inst_cellmath__37_0_I2715 (.Y(inst_cellmath__37[27]), .A0(N3890), .A1(N3966), .B0(N3842), .B1(N3973));
NAND2X1 inst_cellmath__39__19__2mx_I3142 (.Y(N8208), .A(N4277), .B(inst_cellmath__37[27]));
CLKXOR2X1 inst_cellmath__36__15__I7892 (.Y(N13350), .A(N4400), .B(N8208));
INVXL inst_cellmath__36__15__I7893 (.Y(N13359), .A(N13350));
INVXL inst_cellmath__36__15__I7894 (.Y(N13380), .A(N13366));
NOR2XL inst_cellmath__36__15__I7895 (.Y(N13354), .A(N13366), .B(N13350));
NAND2X1 inst_cellmath__36__15__I7896 (.Y(N13365), .A(N13350), .B(N13380));
OR2XL inst_cellmath__36__15__I8135 (.Y(N13372), .A(N13380), .B(N13350));
XOR2XL inst_cellmath__36__15__I7899 (.Y(N4621), .A(N13380), .B(N13359));
INVXL inst_cellmath__36__15__I7900 (.Y(N13385), .A(N4400));
NAND2XL inst_cellmath__37_0_I832 (.Y(N3844), .A(N3977), .B(N3920));
AOI22XL inst_cellmath__37_0_I876 (.Y(inst_cellmath__37[28]), .A0(N3842), .A1(N4022), .B0(N3844), .B1(N3890));
AND2XL inst_cellmath__36__15__I8136 (.Y(N13371), .A(inst_cellmath__37[28]), .B(N4277));
XOR2XL inst_cellmath__36__15__I7903 (.Y(N13369), .A(N13371), .B(N13385));
OR2X1 inst_cellmath__36__15__I7904 (.Y(N13392), .A(N13376), .B(N13369));
XNOR2X1 inst_cellmath__36__15__I7905 (.Y(N13367), .A(N13385), .B(N13371));
XOR2XL inst_cellmath__36__15__I7906 (.Y(N4684), .A(N13384), .B(N13367));
NAND2X2 inst_cellmath__36__15__I7907 (.Y(N13389), .A(N13388), .B(N13375));
INVXL buf1_A_I8282 (.Y(N13872), .A(N13388));
INVXL buf1_A_I8283 (.Y(N4707), .A(N13872));
INVXL buf1_A_I8284 (.Y(N13877), .A(N13375));
INVXL buf1_A_I8285 (.Y(N4639), .A(N13877));
OAI2BB1XL inst_cellmath__36__15__I7910 (.Y(N4657), .A0N(N4707), .A1N(N4639), .B0(N13352));
AOI22X4 inst_cellmath__36__15__I7911 (.Y(N13378), .A0(N13372), .A1(N13365), .B0(N13352), .B1(N13389));
INVXL inst_cellmath__36__15__I7912 (.Y(N13362), .A(N13378));
OAI2BB1X1 inst_cellmath__36__15__I7913 (.Y(N4706), .A0N(N13380), .A1N(N13359), .B0(N13362));
OAI21X4 inst_cellmath__36__15__I7914 (.Y(N13387), .A0(N13354), .A1(N13378), .B0(N4684));
NAND2XL inst_cellmath__37_0_I835 (.Y(N3914), .A(N3920), .B(N3906));
AOI22XL inst_cellmath__37_0_I879 (.Y(inst_cellmath__37[31]), .A0(N3842), .A1(N3945), .B0(N3914), .B1(N3890));
INVXL inst_cellmath__36__15__I8033 (.Y(N13149), .A(N13145));
MXI2XL inst_cellmath__36__15__I8034 (.Y(N13613), .A(a_man[4]), .B(b_man[4]), .S0(N13149));
NAND2XL inst_cellmath__37_0_I834 (.Y(N4034), .A(N3920), .B(N3857));
AOI22XL inst_cellmath__37_0_I878 (.Y(inst_cellmath__37[30]), .A0(N3842), .A1(N3902), .B0(N4034), .B1(N3890));
NAND2XL inst_cellmath__33_49_24_I905 (.Y(inst_cellmath__33[30]), .A(N4277), .B(inst_cellmath__37[30]));
XNOR2X1 inst_cellmath__36__15__I8037 (.Y(N13634), .A(N4400), .B(inst_cellmath__33[30]));
AND2XL inst_cellmath__36__15__I8137 (.Y(N13617), .A(N4277), .B(inst_cellmath__37[31]));
INVXL inst_cellmath__36__15__I8039 (.Y(N13597), .A(N4400));
OR2XL inst_cellmath__36__15__I8190 (.Y(N13615), .A(N13597), .B(N13617));
NAND2XL inst_cellmath__36__15__I8043 (.Y(N13607), .A(N13597), .B(N13617));
XOR2XL inst_cellmath__36__15__I8044 (.Y(N13593), .A(N13597), .B(N13617));
MXI2XL cynw_cm_float_add2_ieee_I952 (.Y(N658), .A(a_man[3]), .B(b_man[3]), .S0(N13149));
NAND2XL inst_cellmath__37_0_I833 (.Y(N3940), .A(N3920), .B(N4026));
AOI22XL inst_cellmath__37_0_I877 (.Y(inst_cellmath__37[29]), .A0(N3842), .A1(N3853), .B0(N3940), .B1(N3890));
NAND2XL inst_cellmath__33_49_24_I904 (.Y(inst_cellmath__33[29]), .A(N4277), .B(inst_cellmath__37[29]));
XNOR2X1 inst_cellmath__39__19__2mx_I977 (.Y(inst_cellmath__39[4]), .A(inst_cellmath__33[29]), .B(N4400));
NAND2XL inst_cellmath__36__15__I8045 (.Y(N13604), .A(N658), .B(inst_cellmath__39[4]));
CLKXOR2X2 inst_cellmath__36__15__I8046 (.Y(N4604), .A(inst_cellmath__39[4]), .B(N658));
AND2XL inst_cellmath__36__15__I8047 (.Y(N13596), .A(N13613), .B(N13634));
XOR2XL inst_cellmath__36__15__I8048 (.Y(N4668), .A(N13613), .B(N13634));
MX2XL inst_cellmath__36__15__I8191 (.Y(N13629), .A(a_man[5]), .B(b_man[5]), .S0(N13149));
AOI21X2 inst_cellmath__36__15__I8052 (.Y(N13621), .A0(N13607), .A1(N13615), .B0(N13629));
XOR2XL inst_cellmath__36__15__I8053 (.Y(N4586), .A(N13629), .B(N13593));
NAND2X4 inst_cellmath__36__15__I8054 (.Y(N13599), .A(N13392), .B(N13387));
INVX2 inst_cellmath__36__15__I8055 (.Y(N13608), .A(N13604));
AOI21X4 inst_cellmath__36__15__I8056 (.Y(N13610), .A0(N4604), .A1(N13599), .B0(N13608));
DLY1X1 inst_cellmath__36__15__I8057 (.Y(N4667), .A(N13599));
OAI2BB1X1 inst_cellmath__36__15__I8058 (.Y(N4691), .A0N(N4604), .A1N(N4667), .B0(N13604));
NOR2BX2 inst_cellmath__36__15__I8059 (.Y(N13627), .AN(N4668), .B(N13610));
INVXL inst_cellmath__36__15__I8060 (.Y(N13611), .A(N13627));
NOR2X2 inst_cellmath__36__15__I8061 (.Y(N13635), .A(N13596), .B(N13627));
OAI2BB1X1 inst_cellmath__36__15__I8062 (.Y(N4635), .A0N(N13613), .A1N(N13634), .B0(N13611));
NOR2BX2 inst_cellmath__36__15__I8063 (.Y(N13601), .AN(N4586), .B(N13635));
NOR2X2 inst_cellmath__36__15__I8064 (.Y(N13606), .A(N13621), .B(N13601));
CLKINVX1 inst_cellmath__36__15__I8065 (.Y(N4643), .A(N13606));
INVXL inst_cellmath__36__15__I7658 (.Y(N13148), .A(N13145));
INVXL inst_cellmath__36__15__I7657 (.Y(N13147), .A(N13145));
INVXL inst_cellmath__36__15__I7656 (.Y(N13146), .A(N13145));
NAND2XL inst_cellmath__37_0_I836 (.Y(N4007), .A(N3949), .B(N3920));
NAND2XL inst_cellmath__37_0_I837 (.Y(N3885), .A(N3920), .B(N3998));
NAND2XL inst_cellmath__37_0_I838 (.Y(N3978), .A(N3920), .B(N4046));
NAND2XL inst_cellmath__37_0_I839 (.Y(N3859), .A(N3876), .B(N3920));
NAND2XL inst_cellmath__37_0_I840 (.Y(N3951), .A(N3925), .B(N3920));
NAND2XL inst_cellmath__37_0_I841 (.Y(N4048), .A(N3920), .B(N3970));
NAND2XL inst_cellmath__37_0_I842 (.Y(N3927), .A(N4016), .B(N3920));
NAND2XL inst_cellmath__37_0_I843 (.Y(N4018), .A(N3848), .B(N3920));
NAND2XL inst_cellmath__37_0_I844 (.Y(N3897), .A(N3895), .B(N3920));
NAND2XL inst_cellmath__37_0_I845 (.Y(N3988), .A(N4037), .B(N3920));
AOI22XL inst_cellmath__37_0_I880 (.Y(inst_cellmath__37[32]), .A0(N3842), .A1(N3994), .B0(N4007), .B1(N3890));
AOI22XL inst_cellmath__37_0_I881 (.Y(inst_cellmath__37[33]), .A0(N3842), .A1(N4042), .B0(N3885), .B1(N3890));
AOI22XL inst_cellmath__37_0_I882 (.Y(inst_cellmath__37[34]), .A0(N3842), .A1(N3872), .B0(N3978), .B1(N3890));
AOI22XL inst_cellmath__37_0_I883 (.Y(inst_cellmath__37[35]), .A0(N3842), .A1(N3966), .B0(N3859), .B1(N3890));
AOI22XL inst_cellmath__37_0_I884 (.Y(inst_cellmath__37[36]), .A0(N3842), .A1(N3844), .B0(N3951), .B1(N3890));
AOI22XL inst_cellmath__37_0_I885 (.Y(inst_cellmath__37[37]), .A0(N3842), .A1(N3940), .B0(N4048), .B1(N3890));
AOI22XL inst_cellmath__37_0_I886 (.Y(inst_cellmath__37[38]), .A0(N3842), .A1(N4034), .B0(N3927), .B1(N3890));
AOI22XL inst_cellmath__37_0_I887 (.Y(inst_cellmath__37[39]), .A0(N3842), .A1(N3914), .B0(N4018), .B1(N3890));
AOI22XL inst_cellmath__37_0_I888 (.Y(inst_cellmath__37[40]), .A0(N3842), .A1(N4007), .B0(N3897), .B1(N3890));
AOI22XL inst_cellmath__37_0_I889 (.Y(inst_cellmath__37[41]), .A0(N3842), .A1(N3885), .B0(N3988), .B1(N3890));
NOR2XL inst_cellmath__37_0_I891 (.Y(inst_cellmath__37[43]), .A(N3890), .B(N3859));
NOR2XL inst_cellmath__37_0_I892 (.Y(inst_cellmath__37[44]), .A(N3890), .B(N3951));
NAND2XL inst_cellmath__33_49_24_I909 (.Y(inst_cellmath__33[34]), .A(N4277), .B(inst_cellmath__37[34]));
NAND2XL inst_cellmath__33_49_24_I910 (.Y(inst_cellmath__33[35]), .A(N4277), .B(inst_cellmath__37[35]));
NAND2XL inst_cellmath__33_49_24_I913 (.Y(inst_cellmath__33[38]), .A(N4277), .B(inst_cellmath__37[38]));
NAND2XL inst_cellmath__33_49_24_I914 (.Y(inst_cellmath__33[39]), .A(N4277), .B(inst_cellmath__37[39]));
NAND2XL inst_cellmath__33_49_24_I915 (.Y(inst_cellmath__33[40]), .A(N4277), .B(inst_cellmath__37[40]));
NOR3BXL inst_cellmath__33_49_24_I2974 (.Y(inst_cellmath__33[42]), .AN(N4277), .B(N3890), .C(N3978));
NAND2XL inst_cellmath__33_49_24_I918 (.Y(inst_cellmath__33[43]), .A(N4277), .B(inst_cellmath__37[43]));
NAND2XL inst_cellmath__33_49_24_I919 (.Y(inst_cellmath__33[44]), .A(N4277), .B(inst_cellmath__37[44]));
NOR3BXL inst_cellmath__33_49_24_I2975 (.Y(inst_cellmath__33[45]), .AN(N4277), .B(N3890), .C(N4048));
NOR3BXL inst_cellmath__33_49_24_I2976 (.Y(inst_cellmath__33[46]), .AN(N4277), .B(N3890), .C(N3927));
NOR3BXL inst_cellmath__33_49_24_I2977 (.Y(inst_cellmath__33[47]), .AN(N4277), .B(N3890), .C(N4018));
NOR3BXL inst_cellmath__33_49_24_I2978 (.Y(inst_cellmath__33[48]), .AN(N4277), .B(N3890), .C(N3897));
NOR3BXL inst_cellmath__33_49_24_I2979 (.Y(inst_cellmath__33[49]), .AN(N4277), .B(N3890), .C(N3988));
MX2XL cynw_cm_float_add2_ieee_I955 (.Y(N661), .A(a_man[6]), .B(b_man[6]), .S0(N13149));
MX2XL cynw_cm_float_add2_ieee_I956 (.Y(N662), .A(a_man[7]), .B(b_man[7]), .S0(N13149));
MXI2XL cynw_cm_float_add2_ieee_I957 (.Y(N663), .A(a_man[8]), .B(b_man[8]), .S0(N13148));
MXI2XL cynw_cm_float_add2_ieee_I958 (.Y(N664), .A(a_man[9]), .B(b_man[9]), .S0(N13148));
MX2XL cynw_cm_float_add2_ieee_I959 (.Y(N665), .A(a_man[10]), .B(b_man[10]), .S0(N13148));
MX2XL cynw_cm_float_add2_ieee_I960 (.Y(N666), .A(a_man[11]), .B(b_man[11]), .S0(N13148));
MXI2XL cynw_cm_float_add2_ieee_I961 (.Y(N667), .A(a_man[12]), .B(b_man[12]), .S0(N13148));
MXI2XL cynw_cm_float_add2_ieee_I962 (.Y(N668), .A(a_man[13]), .B(b_man[13]), .S0(N13147));
MXI2XL cynw_cm_float_add2_ieee_I963 (.Y(N669), .A(a_man[14]), .B(b_man[14]), .S0(N13147));
MX2XL cynw_cm_float_add2_ieee_I964 (.Y(N670), .A(a_man[15]), .B(b_man[15]), .S0(N13147));
MX2XL cynw_cm_float_add2_ieee_I965 (.Y(N671), .A(a_man[16]), .B(b_man[16]), .S0(N13147));
MXI2XL cynw_cm_float_add2_ieee_I966 (.Y(N672), .A(a_man[17]), .B(b_man[17]), .S0(N13147));
MXI2XL cynw_cm_float_add2_ieee_I967 (.Y(N673), .A(a_man[18]), .B(b_man[18]), .S0(N13146));
MX2XL cynw_cm_float_add2_ieee_I968 (.Y(N674), .A(a_man[19]), .B(b_man[19]), .S0(N13146));
MX2XL cynw_cm_float_add2_ieee_I969 (.Y(N675), .A(a_man[20]), .B(b_man[20]), .S0(N13146));
MX2XL cynw_cm_float_add2_ieee_I970 (.Y(N676), .A(a_man[21]), .B(b_man[21]), .S0(N13146));
MX2XL cynw_cm_float_add2_ieee_I971 (.Y(N677), .A(a_man[22]), .B(b_man[22]), .S0(N13146));
NAND2XL node_cs_const1_cs_ii_A_I3146 (.Y(N8222), .A(N4277), .B(inst_cellmath__37[32]));
XOR2XL node_cs_const1_cs_ii_A_I3147 (.Y(inst_cellmath__39[7]), .A(N4400), .B(N8222));
NAND2XL node_cs_const1_cs_ii_A_I3148 (.Y(N8229), .A(N4277), .B(inst_cellmath__37[33]));
XOR2XL node_cs_const1_cs_ii_A_I3149 (.Y(inst_cellmath__39[8]), .A(N4400), .B(N8229));
XNOR2X1 inst_cellmath__39__19__2mx_I982 (.Y(inst_cellmath__39[9]), .A(inst_cellmath__33[34]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I983 (.Y(inst_cellmath__39[10]), .A(inst_cellmath__33[35]), .B(N4400));
NAND2XL node_cs_const1_cs_ii_A_I3150 (.Y(N8236), .A(N4277), .B(inst_cellmath__37[36]));
XOR2XL node_cs_const1_cs_ii_A_I3151 (.Y(inst_cellmath__39[11]), .A(N4400), .B(N8236));
NAND2XL node_cs_const1_cs_ii_A_I3152 (.Y(N8243), .A(N4277), .B(inst_cellmath__37[37]));
XOR2XL node_cs_const1_cs_ii_A_I3153 (.Y(inst_cellmath__39[12]), .A(N4400), .B(N8243));
XNOR2X1 inst_cellmath__39__19__2mx_I986 (.Y(inst_cellmath__39[13]), .A(inst_cellmath__33[38]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I987 (.Y(inst_cellmath__39[14]), .A(inst_cellmath__33[39]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I988 (.Y(inst_cellmath__39[15]), .A(inst_cellmath__33[40]), .B(N4400));
NAND2XL node_cs_const1_cs_ii_A_I3154 (.Y(N8250), .A(N4277), .B(inst_cellmath__37[41]));
XOR2XL node_cs_const1_cs_ii_A_I3155 (.Y(inst_cellmath__39[16]), .A(N4400), .B(N8250));
XNOR2X1 inst_cellmath__39__19__2mx_I990 (.Y(inst_cellmath__39[17]), .A(inst_cellmath__33[42]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I991 (.Y(inst_cellmath__39[18]), .A(inst_cellmath__33[43]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I992 (.Y(inst_cellmath__39[19]), .A(inst_cellmath__33[44]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I993 (.Y(inst_cellmath__39[20]), .A(inst_cellmath__33[45]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I994 (.Y(inst_cellmath__39[21]), .A(inst_cellmath__33[46]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I995 (.Y(inst_cellmath__39[22]), .A(inst_cellmath__33[47]), .B(N4400));
XNOR2X1 inst_cellmath__39__19__2mx_I996 (.Y(inst_cellmath__39[23]), .A(inst_cellmath__33[48]), .B(N4400));
OR2XL inst_cellmath__45_0_I1011 (.Y(N4719), .A(N661), .B(inst_cellmath__39[7]));
XOR2XL inst_cellmath__45_0_I1012 (.Y(N4648), .A(N661), .B(inst_cellmath__39[7]));
OR2XL inst_cellmath__45_0_I1013 (.Y(N4647), .A(N662), .B(inst_cellmath__39[8]));
XOR2XL inst_cellmath__45_0_I1014 (.Y(N4713), .A(N662), .B(inst_cellmath__39[8]));
NAND2XL inst_cellmath__45_0_I1015 (.Y(N4579), .A(N663), .B(inst_cellmath__39[9]));
XOR2XL inst_cellmath__45_0_I1016 (.Y(N4628), .A(N663), .B(inst_cellmath__39[9]));
NAND2XL inst_cellmath__45_0_I1017 (.Y(N4653), .A(N664), .B(inst_cellmath__39[10]));
XOR2XL inst_cellmath__45_0_I1018 (.Y(N4692), .A(N664), .B(inst_cellmath__39[10]));
OR2XL inst_cellmath__45_0_I1019 (.Y(N4589), .A(N665), .B(inst_cellmath__39[11]));
XOR2XL inst_cellmath__45_0_I1020 (.Y(N4610), .A(N665), .B(inst_cellmath__39[11]));
OR2XL inst_cellmath__45_0_I1021 (.Y(N4663), .A(N666), .B(inst_cellmath__39[12]));
XOR2XL inst_cellmath__45_0_I1022 (.Y(N4676), .A(N666), .B(inst_cellmath__39[12]));
NAND2XL inst_cellmath__45_0_I1023 (.Y(N4595), .A(N667), .B(inst_cellmath__39[13]));
XOR2XL inst_cellmath__45_0_I1024 (.Y(N4593), .A(N667), .B(inst_cellmath__39[13]));
NAND2XL inst_cellmath__45_0_I1025 (.Y(N4673), .A(N668), .B(inst_cellmath__39[14]));
XOR2XL inst_cellmath__45_0_I1026 (.Y(N4654), .A(N668), .B(inst_cellmath__39[14]));
NAND2XL inst_cellmath__45_0_I1027 (.Y(N4603), .A(N669), .B(inst_cellmath__39[15]));
XOR2XL inst_cellmath__45_0_I1028 (.Y(N4722), .A(N669), .B(inst_cellmath__39[15]));
OR2XL inst_cellmath__45_0_I1029 (.Y(N4679), .A(N670), .B(inst_cellmath__39[16]));
XOR2XL inst_cellmath__45_0_I1030 (.Y(N4636), .A(N670), .B(inst_cellmath__39[16]));
OR2XL inst_cellmath__45_0_I1031 (.Y(N4609), .A(N671), .B(inst_cellmath__39[17]));
XOR2XL inst_cellmath__45_0_I1032 (.Y(N4700), .A(N671), .B(inst_cellmath__39[17]));
NAND2XL inst_cellmath__45_0_I1033 (.Y(N4687), .A(N672), .B(inst_cellmath__39[18]));
XOR2XL inst_cellmath__45_0_I1034 (.Y(N4620), .A(N672), .B(inst_cellmath__39[18]));
NAND2XL inst_cellmath__45_0_I1035 (.Y(N4618), .A(N673), .B(inst_cellmath__39[19]));
XOR2XL inst_cellmath__45_0_I1036 (.Y(N4682), .A(N673), .B(inst_cellmath__39[19]));
OR2XL inst_cellmath__45_0_I1037 (.Y(N4695), .A(N674), .B(inst_cellmath__39[20]));
XOR2XL inst_cellmath__45_0_I1038 (.Y(N4600), .A(N674), .B(inst_cellmath__39[20]));
OR2XL inst_cellmath__45_0_I1039 (.Y(N4626), .A(N675), .B(inst_cellmath__39[21]));
XOR2XL inst_cellmath__45_0_I1040 (.Y(N4665), .A(N675), .B(inst_cellmath__39[21]));
OR2XL inst_cellmath__45_0_I1041 (.Y(N4704), .A(N676), .B(inst_cellmath__39[22]));
XOR2XL inst_cellmath__45_0_I1042 (.Y(N4582), .A(N676), .B(inst_cellmath__39[22]));
XOR2XL inst_cellmath__45_0_I1044 (.Y(N4644), .A(N677), .B(inst_cellmath__39[23]));
CLKXOR2X1 inst_cellmath__45_0_I2991 (.Y(N4677), .A(N4400), .B(inst_cellmath__33[49]));
OAI2BB1XL inst_cellmath__45_0_I1052 (.Y(N4718), .A0N(N4648), .A1N(N4643), .B0(N4719));
OAI2BB1XL inst_cellmath__45_0_I1053 (.Y(N4709), .A0N(N4713), .A1N(N4718), .B0(N4647));
OAI2BB1XL inst_cellmath__45_0_I1054 (.Y(N4612), .A0N(N4628), .A1N(N4709), .B0(N4579));
OAI2BB1XL inst_cellmath__45_0_I1055 (.Y(N4583), .A0N(N4692), .A1N(N4612), .B0(N4653));
OAI2BB1XL inst_cellmath__45_0_I1056 (.Y(N4616), .A0N(N4610), .A1N(N4583), .B0(N4589));
OAI2BB1XL inst_cellmath__45_0_I1057 (.Y(N4717), .A0N(N4676), .A1N(N4616), .B0(N4663));
OAI2BB1XL inst_cellmath__45_0_I1058 (.Y(N4585), .A0N(N4593), .A1N(N4717), .B0(N4595));
OAI2BB1XL inst_cellmath__45_0_I1059 (.Y(N4664), .A0N(N4654), .A1N(N4585), .B0(N4673));
OAI2BB1X1 inst_cellmath__45_0_I1060 (.Y(N4659), .A0N(N4722), .A1N(N4664), .B0(N4603));
OAI2BB1X1 inst_cellmath__45_0_I1061 (.Y(N4723), .A0N(N4636), .A1N(N4659), .B0(N4679));
OAI2BB1X1 inst_cellmath__45_0_I1062 (.Y(N4699), .A0N(N4700), .A1N(N4723), .B0(N4609));
OAI2BB1X1 inst_cellmath__45_0_I1063 (.Y(N4597), .A0N(N4620), .A1N(N4699), .B0(N4687));
OAI2BB1X1 inst_cellmath__45_0_I1064 (.Y(N4701), .A0N(N4682), .A1N(N4597), .B0(N4618));
OAI2BB1X1 inst_cellmath__45_0_I1065 (.Y(N4578), .A0N(N4600), .A1N(N4701), .B0(N4695));
OAI2BB1X1 inst_cellmath__45_0_I1066 (.Y(N4666), .A0N(N4665), .A1N(N4578), .B0(N4626));
OAI2BB1X1 inst_cellmath__45_0_I1067 (.Y(N4672), .A0N(N4582), .A1N(N4666), .B0(N4704));
OR2XL gen2_alt_A_I8148 (.Y(N8257), .A(N677), .B(inst_cellmath__39[23]));
OAI2BB1X1 gen2_alt_A_I3157 (.Y(N4594), .A0N(N4644), .A1N(N4672), .B0(N8257));
XOR2XL inst_cellmath__45_0_I1069 (.Y(inst_cellmath__45[0]), .A(inst_cellmath__44), .B(inst_cellmath__39[0]));
XNOR2X1 inst_cellmath__45_0_I1070 (.Y(inst_cellmath__45[1]), .A(N4639), .B(N4707));
XNOR2X1 inst_cellmath__45_0_I1071 (.Y(inst_cellmath__45[2]), .A(N4657), .B(N4621));
XNOR2X1 inst_cellmath__45_0_I1072 (.Y(inst_cellmath__45[3]), .A(N4706), .B(N4684));
XNOR2X1 inst_cellmath__45_0_I1073 (.Y(inst_cellmath__45[4]), .A(N4667), .B(N4604));
XNOR2X1 inst_cellmath__45_0_I1074 (.Y(inst_cellmath__45[5]), .A(N4691), .B(N4668));
XNOR2X1 inst_cellmath__45_0_I1075 (.Y(inst_cellmath__45[6]), .A(N4635), .B(N4586));
XNOR2X1 inst_cellmath__45_0_I1076 (.Y(inst_cellmath__45[7]), .A(N4643), .B(N4648));
XNOR2X1 inst_cellmath__45_0_I1077 (.Y(inst_cellmath__45[8]), .A(N4718), .B(N4713));
XNOR2X1 inst_cellmath__45_0_I1078 (.Y(inst_cellmath__45[9]), .A(N4709), .B(N4628));
XNOR2X1 inst_cellmath__45_0_I1079 (.Y(inst_cellmath__45[10]), .A(N4612), .B(N4692));
XNOR2X1 inst_cellmath__45_0_I1080 (.Y(inst_cellmath__45[11]), .A(N4583), .B(N4610));
XNOR2X1 inst_cellmath__45_0_I1081 (.Y(inst_cellmath__45[12]), .A(N4616), .B(N4676));
XNOR2X1 inst_cellmath__45_0_I1082 (.Y(inst_cellmath__45[13]), .A(N4717), .B(N4593));
XNOR2X1 inst_cellmath__45_0_I1083 (.Y(inst_cellmath__45[14]), .A(N4585), .B(N4654));
XNOR2X1 inst_cellmath__45_0_I1084 (.Y(inst_cellmath__45[15]), .A(N4664), .B(N4722));
XNOR2X1 inst_cellmath__45_0_I1085 (.Y(inst_cellmath__45[16]), .A(N4659), .B(N4636));
XNOR2X1 inst_cellmath__45_0_I1086 (.Y(inst_cellmath__45[17]), .A(N4723), .B(N4700));
XNOR2X1 inst_cellmath__45_0_I1087 (.Y(inst_cellmath__45[18]), .A(N4699), .B(N4620));
XNOR2X1 inst_cellmath__45_0_I1088 (.Y(inst_cellmath__45[19]), .A(N4597), .B(N4682));
XNOR2X1 inst_cellmath__45_0_I1089 (.Y(inst_cellmath__45[20]), .A(N4701), .B(N4600));
XNOR2X1 inst_cellmath__45_0_I1090 (.Y(inst_cellmath__45[21]), .A(N4578), .B(N4665));
XNOR2XL inst_cellmath__45_0_I1091 (.Y(inst_cellmath__45[22]), .A(N4666), .B(N4582));
XNOR2X1 inst_cellmath__45_0_I1092 (.Y(inst_cellmath__45[23]), .A(N4672), .B(N4644));
XNOR2X1 inst_cellmath__45_0_I1093 (.Y(inst_cellmath__45[24]), .A(N4594), .B(N4677));
NAND2X1 inst_cellmath__45_0_I1094 (.Y(N4624), .A(N4677), .B(N4594));
CLKXOR2X1 inst_cellmath__45_0_I1095 (.Y(inst_cellmath__45[25]), .A(inst_cellmath__39[25]), .B(N4624));
NOR2BX1 inst_cellmath__49_0_I1096 (.Y(N4848), .AN(inst_cellmath__45[0]), .B(inst_cellmath__45[1]));
NOR2XL inst_cellmath__49_0_I1097 (.Y(N4827), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[0]));
NOR2BX1 inst_cellmath__49_0_I1098 (.Y(N4869), .AN(inst_cellmath__45[2]), .B(inst_cellmath__45[3]));
INVXL inst_cellmath__49_0_I1099 (.Y(N4888), .A(inst_cellmath__45[5]));
OAI21XL inst_cellmath__49_0_I1100 (.Y(N4910), .A0(inst_cellmath__45[4]), .A1(N4869), .B0(N4888));
NOR2XL inst_cellmath__49_0_I1101 (.Y(N4837), .A(inst_cellmath__45[3]), .B(inst_cellmath__45[2]));
NOR2XL inst_cellmath__49_0_I1102 (.Y(N4856), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[4]));
NOR2BX1 inst_cellmath__49_0_I1103 (.Y(N4898), .AN(inst_cellmath__45[6]), .B(inst_cellmath__45[7]));
INVXL inst_cellmath__49_0_I1104 (.Y(N4918), .A(inst_cellmath__45[9]));
OAI21XL inst_cellmath__49_0_I1105 (.Y(N4846), .A0(inst_cellmath__45[8]), .A1(N4898), .B0(N4918));
NOR2XL inst_cellmath__49_0_I1106 (.Y(N4864), .A(inst_cellmath__45[7]), .B(inst_cellmath__45[6]));
NOR2XL inst_cellmath__49_0_I1107 (.Y(N4883), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[8]));
NOR2BX1 inst_cellmath__49_0_I1108 (.Y(N4832), .AN(inst_cellmath__45[10]), .B(inst_cellmath__45[11]));
INVXL inst_cellmath__49_0_I1109 (.Y(N4852), .A(inst_cellmath__45[13]));
OAI21XL inst_cellmath__49_0_I1110 (.Y(N4874), .A0(inst_cellmath__45[12]), .A1(N4832), .B0(N4852));
NOR2XL inst_cellmath__49_0_I1111 (.Y(N4894), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[10]));
NOR2XL inst_cellmath__49_0_I1112 (.Y(N4914), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[12]));
NOR2BX1 inst_cellmath__49_0_I1113 (.Y(N4860), .AN(inst_cellmath__45[14]), .B(inst_cellmath__45[15]));
INVXL inst_cellmath__49_0_I1114 (.Y(N4881), .A(inst_cellmath__45[17]));
OAI21XL inst_cellmath__49_0_I1115 (.Y(N4902), .A0(inst_cellmath__45[16]), .A1(N4860), .B0(N4881));
NOR2XL inst_cellmath__49_0_I1116 (.Y(N4829), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[14]));
NOR2XL inst_cellmath__49_0_I1117 (.Y(N4850), .A(inst_cellmath__45[17]), .B(inst_cellmath__45[16]));
NOR2BX1 inst_cellmath__49_0_I1118 (.Y(N4889), .AN(inst_cellmath__45[18]), .B(inst_cellmath__45[19]));
INVXL inst_cellmath__49_0_I1119 (.Y(N4911), .A(inst_cellmath__45[21]));
OAI21XL inst_cellmath__49_0_I1120 (.Y(N4838), .A0(inst_cellmath__45[20]), .A1(N4889), .B0(N4911));
NOR2XL inst_cellmath__49_0_I1121 (.Y(N4857), .A(inst_cellmath__45[19]), .B(inst_cellmath__45[18]));
NOR2XL inst_cellmath__49_0_I1122 (.Y(N4878), .A(inst_cellmath__45[21]), .B(inst_cellmath__45[20]));
NOR2BX1 inst_cellmath__49_0_I1123 (.Y(N4824), .AN(inst_cellmath__45[22]), .B(inst_cellmath__45[23]));
INVXL inst_cellmath__49_0_I1124 (.Y(N4847), .A(inst_cellmath__45[25]));
OAI21X1 inst_cellmath__49_0_I1125 (.Y(N4866), .A0(N4824), .A1(inst_cellmath__45[24]), .B0(N4847));
NOR2X4 inst_cellmath__49_0_I1126 (.Y(N4885), .A(inst_cellmath__45[23]), .B(inst_cellmath__45[22]));
NOR2X2 inst_cellmath__49_0_I1127 (.Y(N4907), .A(inst_cellmath__45[25]), .B(inst_cellmath__45[24]));
NAND2BXL inst_cellmath__49_0_I1128 (.Y(N4904), .AN(N4837), .B(N4856));
NAND2XL inst_cellmath__49_0_I1129 (.Y(N4872), .A(N4856), .B(N4837));
NAND2XL inst_cellmath__49_0_I1130 (.Y(N4891), .A(N4883), .B(N4864));
NAND2BXL inst_cellmath__49_0_I1131 (.Y(N4840), .AN(N4894), .B(N4914));
INVXL inst_cellmath__49_0_I1132 (.Y(N4859), .A(N4850));
AOI21XL inst_cellmath__49_0_I1133 (.Y(N4880), .A0(N4829), .A1(N4840), .B0(N4859));
NAND2XL inst_cellmath__49_0_I1134 (.Y(N4900), .A(N4914), .B(N4894));
NAND2XL inst_cellmath__49_0_I1135 (.Y(N4826), .A(N4850), .B(N4829));
NAND2BXL inst_cellmath__49_0_I1136 (.Y(N4868), .AN(N4857), .B(N4878));
INVXL inst_cellmath__49_0_I1137 (.Y(N4887), .A(N4907));
AOI21XL inst_cellmath__49_0_I1138 (.Y(N4909), .A0(N4885), .A1(N4868), .B0(N4887));
NAND2X4 inst_cellmath__49_0_I1139 (.Y(N4836), .A(N4878), .B(N4857));
NAND2X4 inst_cellmath__49_0_I1140 (.Y(N4855), .A(N4885), .B(N4907));
NAND2BXL inst_cellmath__49_0_I1141 (.Y(N4845), .AN(N4891), .B(N4872));
NOR2XL inst_cellmath__49_0_I1142 (.Y(N4831), .A(N4891), .B(N4872));
NOR2BX1 inst_cellmath__49_0_I1143 (.Y(N4873), .AN(N4900), .B(N4826));
INVXL inst_cellmath__49_0_I1144 (.Y(N4893), .A(N4855));
OAI21XL inst_cellmath__49_0_I1145 (.Y(N4913), .A0(N4836), .A1(N4873), .B0(N4893));
NOR2X2 inst_cellmath__49_0_I1146 (.Y(N4842), .A(N4826), .B(N4900));
NOR2X6 inst_cellmath__49_0_I1147 (.Y(N4892), .A(N4836), .B(N4855));
NAND2BXL inst_cellmath__49_0_I1148 (.Y(N4901), .AN(N4827), .B(N4831));
INVX1 inst_cellmath__49_0_I1149 (.Y(N4828), .A(N4892));
OAI2BB1X1 inst_cellmath__49_0_I1156 (.Y(N4896), .A0N(N4864), .A1N(N4904), .B0(N4883));
AOI21XL inst_cellmath__49_0_I1157 (.Y(N4862), .A0(N4892), .A1(N4880), .B0(N4909));
OAI21XL inst_cellmath__49_0_I1159 (.Y(N4835), .A0(N4891), .A1(N4910), .B0(N4846));
OAI21XL inst_cellmath__49_0_I1160 (.Y(N4877), .A0(N4826), .A1(N4874), .B0(N4902));
OAI21X1 inst_cellmath__49_0_I1161 (.Y(N4917), .A0(N4838), .A1(N4855), .B0(N4866));
AOI21XL inst_cellmath__49_0_I1162 (.Y(N4863), .A0(N4831), .A1(N4848), .B0(N4835));
AOI21X2 inst_cellmath__49_0_I1163 (.Y(N4905), .A0(N4877), .A1(N4892), .B0(N4917));
NAND2X4 inst_cellmath__59_0_I8072 (.Y(N4841), .A(N4842), .B(N4892));
OAI21X2 inst_cellmath__49_0_I1164 (.Y(inst_cellmath__49[0]), .A0(N4863), .A1(N4841), .B0(N4905));
NAND2X1 inst_cellmath__59_0_I8071 (.Y(N4870), .A(N4827), .B(N4831));
NOR2XL inst_cellmath__59_0_I8073 (.Y(inst_cellmath__49[5]), .A(N4870), .B(N4841));
OR2XL cmp_A_I8286 (.Y(N13881), .A(a_sign), .B(b_sign));
AO22XL cmp_A_I8287 (.Y(N645), .A0(N13881), .A1(inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL cynw_cm_float_add2_ieee_I1170 (.Y(inst_cellmath__66), .A(inst_cellmath__11), .B(inst_cellmath__16), .C(N645));
NOR2BX1 inst_cellmath__64__48__2WWMM_I1171 (.Y(N5043), .AN(inst_cellmath__18), .B(inst_cellmath__13));
AOI22XL inst_cellmath__64__48__2WWMM_I1172 (.Y(N5064), .A0(a_sign), .A1(inst_cellmath__13), .B0(N5043), .B1(b_sign));
AO22XL inst_cellmath__64__48__2WWMM_I1173 (.Y(inst_cellmath__64[0]), .A0(inst_cellmath__13), .A1(a_man[0]), .B0(N5043), .B1(b_man[0]));
AO22XL inst_cellmath__64__48__2WWMM_I1174 (.Y(inst_cellmath__64[1]), .A0(inst_cellmath__13), .A1(a_man[1]), .B0(N5043), .B1(b_man[1]));
AO22XL inst_cellmath__64__48__2WWMM_I1175 (.Y(inst_cellmath__64[2]), .A0(inst_cellmath__13), .A1(a_man[2]), .B0(N5043), .B1(b_man[2]));
AO22XL inst_cellmath__64__48__2WWMM_I1176 (.Y(inst_cellmath__64[3]), .A0(inst_cellmath__13), .A1(a_man[3]), .B0(N5043), .B1(b_man[3]));
AO22XL inst_cellmath__64__48__2WWMM_I1177 (.Y(inst_cellmath__64[4]), .A0(inst_cellmath__13), .A1(a_man[4]), .B0(N5043), .B1(b_man[4]));
AO22XL inst_cellmath__64__48__2WWMM_I1178 (.Y(inst_cellmath__64[5]), .A0(inst_cellmath__13), .A1(a_man[5]), .B0(N5043), .B1(b_man[5]));
AO22XL inst_cellmath__64__48__2WWMM_I1179 (.Y(inst_cellmath__64[6]), .A0(inst_cellmath__13), .A1(a_man[6]), .B0(N5043), .B1(b_man[6]));
AO22XL inst_cellmath__64__48__2WWMM_I1180 (.Y(inst_cellmath__64[7]), .A0(inst_cellmath__13), .A1(a_man[7]), .B0(N5043), .B1(b_man[7]));
AO22XL inst_cellmath__64__48__2WWMM_I1181 (.Y(inst_cellmath__64[8]), .A0(inst_cellmath__13), .A1(a_man[8]), .B0(N5043), .B1(b_man[8]));
AO22XL inst_cellmath__64__48__2WWMM_I1182 (.Y(inst_cellmath__64[9]), .A0(inst_cellmath__13), .A1(a_man[9]), .B0(N5043), .B1(b_man[9]));
AO22XL inst_cellmath__64__48__2WWMM_I1183 (.Y(inst_cellmath__64[10]), .A0(inst_cellmath__13), .A1(a_man[10]), .B0(N5043), .B1(b_man[10]));
AO22XL inst_cellmath__64__48__2WWMM_I1184 (.Y(inst_cellmath__64[11]), .A0(inst_cellmath__13), .A1(a_man[11]), .B0(N5043), .B1(b_man[11]));
AO22XL inst_cellmath__64__48__2WWMM_I1185 (.Y(inst_cellmath__64[12]), .A0(inst_cellmath__13), .A1(a_man[12]), .B0(N5043), .B1(b_man[12]));
AO22XL inst_cellmath__64__48__2WWMM_I1186 (.Y(inst_cellmath__64[13]), .A0(inst_cellmath__13), .A1(a_man[13]), .B0(N5043), .B1(b_man[13]));
AO22XL inst_cellmath__64__48__2WWMM_I1187 (.Y(inst_cellmath__64[14]), .A0(inst_cellmath__13), .A1(a_man[14]), .B0(N5043), .B1(b_man[14]));
AO22XL inst_cellmath__64__48__2WWMM_I1188 (.Y(inst_cellmath__64[15]), .A0(inst_cellmath__13), .A1(a_man[15]), .B0(N5043), .B1(b_man[15]));
AO22XL inst_cellmath__64__48__2WWMM_I1189 (.Y(inst_cellmath__64[16]), .A0(inst_cellmath__13), .A1(a_man[16]), .B0(N5043), .B1(b_man[16]));
AO22XL inst_cellmath__64__48__2WWMM_I1190 (.Y(inst_cellmath__64[17]), .A0(inst_cellmath__13), .A1(a_man[17]), .B0(N5043), .B1(b_man[17]));
AO22XL inst_cellmath__64__48__2WWMM_I1191 (.Y(inst_cellmath__64[18]), .A0(inst_cellmath__13), .A1(a_man[18]), .B0(N5043), .B1(b_man[18]));
AO22XL inst_cellmath__64__48__2WWMM_I1192 (.Y(inst_cellmath__64[19]), .A0(inst_cellmath__13), .A1(a_man[19]), .B0(N5043), .B1(b_man[19]));
AO22XL inst_cellmath__64__48__2WWMM_I1193 (.Y(inst_cellmath__64[20]), .A0(inst_cellmath__13), .A1(a_man[20]), .B0(N5043), .B1(b_man[20]));
AO22XL inst_cellmath__64__48__2WWMM_I1194 (.Y(inst_cellmath__64[21]), .A0(inst_cellmath__13), .A1(a_man[21]), .B0(N5043), .B1(b_man[21]));
OAI21XL inst_cellmath__64__48__2WWMM_I1195 (.Y(N710), .A0(inst_cellmath__18), .A1(inst_cellmath__13), .B0(N5064));
OR3X1 inst_cellmath__59_0_I8069 (.Y(inst_cellmath__63), .A(inst_cellmath__13), .B(inst_cellmath__18), .C(N547));
MX2XL inst_cellmath__67_0_I1196 (.Y(N5113), .A(inst_cellmath__66), .B(N710), .S0(inst_cellmath__63));
AND2XL inst_cellmath__59_0_I8070 (.Y(N706), .A(inst_cellmath__11), .B(inst_cellmath__16));
NOR2XL inst_cellmath__67_0_I1197 (.Y(N5122), .A(inst_cellmath__63), .B(N706));
MX2XL inst_cellmath__67_0_I8150 (.Y(N5116), .A(inst_cellmath__48), .B(inst_cellmath__6), .S0(inst_cellmath__49[5]));
MX2XL inst_cellmath__67_0_I1199 (.Y(x[31]), .A(N5113), .B(N5116), .S0(N5122));
AO21X4 inst_cellmath__50_0_I3100 (.Y(N5270), .A0(N4901), .A1(N4842), .B0(N4828));
CLKINVX4 inst_cellmath__50_0_I2910 (.Y(N8174), .A(N5270));
INVX2 inst_cellmath__50_0_I2916 (.Y(N8180), .A(N8174));
INVX1 inst_cellmath__50_0_I2915 (.Y(N8179), .A(N8174));
INVX1 inst_cellmath__50_0_I2914 (.Y(N8178), .A(N8174));
INVX1 inst_cellmath__50_0_I2913 (.Y(N8177), .A(N8174));
CLKAND2X3 inst_cellmath__50_0_I1201 (.Y(N5143), .A(inst_cellmath__45[0]), .B(N5270));
CLKAND2X2 inst_cellmath__50_0_I1202 (.Y(N5214), .A(inst_cellmath__45[1]), .B(N8180));
CLKAND2X3 inst_cellmath__50_0_I1203 (.Y(N5285), .A(inst_cellmath__45[2]), .B(N8180));
AND2XL inst_cellmath__50_0_I1204 (.Y(N5192), .A(N8180), .B(inst_cellmath__45[3]));
AND2XL inst_cellmath__50_0_I1205 (.Y(N5263), .A(N8180), .B(inst_cellmath__45[4]));
AND2XL inst_cellmath__50_0_I1206 (.Y(N5172), .A(N8179), .B(inst_cellmath__45[5]));
AND2XL inst_cellmath__50_0_I1207 (.Y(N5242), .A(N8179), .B(inst_cellmath__45[6]));
AND2XL inst_cellmath__50_0_I1208 (.Y(N5152), .A(N8179), .B(inst_cellmath__45[7]));
MX2XL inst_cellmath__50_0_I1209 (.Y(N5223), .A(inst_cellmath__45[0]), .B(inst_cellmath__45[8]), .S0(N8179));
MX2XL inst_cellmath__50_0_I1210 (.Y(N5258), .A(inst_cellmath__45[1]), .B(inst_cellmath__45[9]), .S0(N8178));
MX2XL inst_cellmath__50_0_I1211 (.Y(N5128), .A(inst_cellmath__45[2]), .B(inst_cellmath__45[10]), .S0(N8178));
MX2XL inst_cellmath__50_0_I1212 (.Y(N5165), .A(inst_cellmath__45[3]), .B(inst_cellmath__45[11]), .S0(N8178));
MX2XL inst_cellmath__50_0_I1213 (.Y(N5202), .A(inst_cellmath__45[4]), .B(inst_cellmath__45[12]), .S0(N8178));
MX2XL inst_cellmath__50_0_I1214 (.Y(N5236), .A(inst_cellmath__45[5]), .B(inst_cellmath__45[13]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1215 (.Y(N5272), .A(inst_cellmath__45[6]), .B(inst_cellmath__45[14]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1216 (.Y(N5146), .A(inst_cellmath__45[7]), .B(inst_cellmath__45[15]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1217 (.Y(N5180), .A(inst_cellmath__45[8]), .B(inst_cellmath__45[16]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1218 (.Y(N5217), .A(inst_cellmath__45[9]), .B(inst_cellmath__45[17]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1219 (.Y(N5251), .A(inst_cellmath__45[10]), .B(inst_cellmath__45[18]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1220 (.Y(N5288), .A(inst_cellmath__45[11]), .B(inst_cellmath__45[19]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1221 (.Y(N5159), .A(inst_cellmath__45[12]), .B(inst_cellmath__45[20]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1222 (.Y(N5196), .A(inst_cellmath__45[13]), .B(inst_cellmath__45[21]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1223 (.Y(N5231), .A(inst_cellmath__45[14]), .B(inst_cellmath__45[22]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1224 (.Y(N5267), .A(inst_cellmath__45[15]), .B(inst_cellmath__45[23]), .S0(N8177));
MX2XL inst_cellmath__50_0_I1225 (.Y(N5138), .A(inst_cellmath__45[16]), .B(inst_cellmath__45[24]), .S0(N8177));
NAND2BX4 inst_cellmath__50_0_I3043 (.Y(N5142), .AN(N4841), .B(N4870));
INVX1 inst_cellmath__50_0_I1227 (.Y(N5178), .A(N5142));
NAND2X4 inst_cellmath__50_0_I1228 (.Y(N5134), .A(N5142), .B(N5143));
NAND2X8 inst_cellmath__50_0_I1229 (.Y(N5208), .A(N5142), .B(N5214));
NAND2X4 inst_cellmath__50_0_I1230 (.Y(N5278), .A(N5142), .B(N5285));
NAND2XL inst_cellmath__50_0_I1231 (.Y(N5186), .A(N5192), .B(N5142));
NAND2XL inst_cellmath__50_0_I1232 (.Y(N5257), .A(N5263), .B(N5142));
NAND2XL inst_cellmath__50_0_I1233 (.Y(N5164), .A(N5172), .B(N5142));
NAND2XL inst_cellmath__50_0_I1234 (.Y(N5235), .A(N5242), .B(N5142));
NAND2XL inst_cellmath__50_0_I1235 (.Y(N5145), .A(N5152), .B(N5142));
NAND2X1 inst_cellmath__50_0_I1236 (.Y(N5216), .A(N5142), .B(N5223));
NAND2X1 inst_cellmath__50_0_I1237 (.Y(N5287), .A(N5142), .B(N5258));
NAND2X1 inst_cellmath__50_0_I1238 (.Y(N5195), .A(N5142), .B(N5128));
NAND2XL inst_cellmath__50_0_I1239 (.Y(N5266), .A(N5165), .B(N5142));
NAND2X1 inst_cellmath__50_0_I1240 (.Y(N5175), .A(N5142), .B(N5202));
NAND2X1 inst_cellmath__50_0_I1241 (.Y(N5245), .A(N5142), .B(N5236));
NAND2X1 inst_cellmath__50_0_I1242 (.Y(N5155), .A(N5142), .B(N5272));
NAND2XL inst_cellmath__50_0_I1243 (.Y(N5226), .A(N5146), .B(N5142));
AOI22XL inst_cellmath__50_0_I1244 (.Y(N5131), .A0(N5178), .A1(N5143), .B0(N5180), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1245 (.Y(N5168), .A0(N5178), .A1(N5214), .B0(N5217), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1246 (.Y(N5205), .A0(N5178), .A1(N5285), .B0(N5251), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1247 (.Y(N5239), .A0(N5178), .A1(N5192), .B0(N5288), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1248 (.Y(N5275), .A0(N5178), .A1(N5263), .B0(N5159), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1249 (.Y(N5149), .A0(N5178), .A1(N5172), .B0(N5196), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1250 (.Y(N5183), .A0(N5178), .A1(N5242), .B0(N5231), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1251 (.Y(N5220), .A0(N5178), .A1(N5152), .B0(N5267), .B1(N5142));
AOI22XL inst_cellmath__50_0_I1252 (.Y(N5254), .A0(N5178), .A1(N5223), .B0(N5138), .B1(N5142));
INVX3 inst_cellmath__50_0_I1253 (.Y(N5247), .A(inst_cellmath__49[0]));
BUFX3 inst_cellmath__50_0_I3102 (.Y(N8182), .A(N5247));
INVX2 inst_cellmath__50_0_I7661 (.Y(N13151), .A(N8182));
CLKINVX4 inst_cellmath__50_0_I7662 (.Y(N13152), .A(N13151));
CLKINVX4 inst_cellmath__50_0_I1254 (.Y(N5283), .A(N5247));
AOI22XL inst_cellmath__50_0_I1260 (.Y(N5174), .A0(N13152), .A1(N5164), .B0(N5257), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1261 (.Y(N5210), .A0(N13152), .A1(N5235), .B0(N5164), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1262 (.Y(N5243), .A0(N13152), .A1(N5145), .B0(N5235), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1263 (.Y(N5279), .A0(N13152), .A1(N5216), .B0(N5145), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1272 (.Y(N5274), .A0(N13152), .A1(N5168), .B0(N5131), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1273 (.Y(N5148), .A0(N13152), .A1(N5205), .B0(N5168), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1274 (.Y(N5181), .A0(N13152), .A1(N5239), .B0(N5205), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1275 (.Y(N5218), .A0(N13152), .A1(N5275), .B0(N5239), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1276 (.Y(N5253), .A0(N13152), .A1(N5149), .B0(N5275), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1277 (.Y(N5290), .A0(N13152), .A1(N5183), .B0(N5149), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1278 (.Y(N5161), .A0(N13152), .A1(N5220), .B0(N5183), .B1(N5283));
AOI22XL inst_cellmath__50_0_I1279 (.Y(N5198), .A0(N13152), .A1(N5254), .B0(N5220), .B1(N5283));
NOR2X6 inst_cellmath__50_0_I7853 (.Y(N13284), .A(N5134), .B(N5283));
AOI22X2 inst_cellmath__50_0_I7854 (.Y(N5193), .A0(N5208), .A1(N13152), .B0(N5134), .B1(N5283));
AOI22X2 inst_cellmath__50_0_I7855 (.Y(N5229), .A0(N5278), .A1(N8182), .B0(N5208), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7856 (.Y(N5265), .A0(N13152), .A1(N5186), .B0(N5278), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7857 (.Y(N5137), .A0(N13152), .A1(N5257), .B0(N5186), .B1(N5283));
OA21X2 inst_cellmath__50_0_I7988 (.Y(N5191), .A0(N4845), .A1(N4841), .B0(N4913));
NAND2X4 inst_cellmath__50_0_I7860 (.Y(N5139), .A(N5191), .B(N13284));
AND2XL inst_cellmath__50_0_I7861 (.Y(N13298), .A(N5191), .B(N5193));
NAND2X1 inst_cellmath__50_0_I7862 (.Y(N5211), .A(N5191), .B(N5193));
NAND2X2 inst_cellmath__50_0_I7863 (.Y(N13272), .A(N5191), .B(N5229));
AND2XL inst_cellmath__50_0_I7864 (.Y(N13294), .A(N5191), .B(N5265));
NAND2XL inst_cellmath__50_0_I7865 (.Y(N5189), .A(N5265), .B(N5191));
INVX2 inst_cellmath__50_0_I7989 (.Y(N5228), .A(N5191));
AOI22XL inst_cellmath__50_0_I7866 (.Y(N5261), .A0(N5228), .A1(N13284), .B0(N5191), .B1(N5137));
AOI22XL inst_cellmath__50_0_I7980 (.Y(N13486), .A0(N13152), .A1(N5287), .B0(N5216), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7981 (.Y(N13504), .A0(N13152), .A1(N5195), .B0(N5287), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7982 (.Y(N13518), .A0(N13152), .A1(N5266), .B0(N5195), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7983 (.Y(N13533), .A0(N13152), .A1(N5175), .B0(N5266), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7984 (.Y(N5129), .A0(N5245), .A1(N13152), .B0(N5175), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7985 (.Y(N5166), .A0(N13152), .A1(N5155), .B0(N5245), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7986 (.Y(N5204), .A0(N13152), .A1(N5226), .B0(N5155), .B1(N5283));
AOI22XL inst_cellmath__50_0_I7987 (.Y(N5238), .A0(N13152), .A1(N5131), .B0(N5226), .B1(N5283));
INVXL buf1_A_I8288 (.Y(N13889), .A(N5191));
INVXL buf1_A_I8289 (.Y(N13475), .A(N13889));
AOI22X1 inst_cellmath__50_0_I7991 (.Y(N13540), .A0(N5174), .A1(N5228), .B0(N13475), .B1(N13486));
AOI22X1 inst_cellmath__50_0_I7992 (.Y(N13483), .A0(N5210), .A1(N5228), .B0(N13475), .B1(N13504));
AOI22X1 inst_cellmath__50_0_I7993 (.Y(N13500), .A0(N5243), .A1(N5228), .B0(N13518), .B1(N13475));
AOI22X1 inst_cellmath__50_0_I7994 (.Y(N13515), .A0(N5228), .A1(N5279), .B0(N13475), .B1(N13533));
INVXL inst_cellmath__50_0_I7995 (.Y(N13535), .A(N5228));
NAND2X1 inst_cellmath__50_0_I7996 (.Y(N13489), .A(N13535), .B(N5129));
NAND2X1 inst_cellmath__50_0_I7998 (.Y(N13499), .A(N13535), .B(N5166));
AOI22X1 inst_cellmath__50_0_I8000 (.Y(N5162), .A0(N13518), .A1(N5228), .B0(N13535), .B1(N5204));
AOI22X1 inst_cellmath__50_0_I8001 (.Y(N5199), .A0(N13533), .A1(N5228), .B0(N13535), .B1(N5238));
OAI21X2 inst_cellmath__50_0_I8002 (.Y(inst_cellmath__49[1]), .A0(N4841), .A1(N4896), .B0(N4862));
INVX1 inst_cellmath__50_0_I8003 (.Y(N13468), .A(inst_cellmath__49[1]));
INVX3 inst_cellmath__50_0_I8004 (.Y(N5171), .A(N13468));
BUFX8 inst_cellmath__50_0_I8005 (.Y(N5135), .A(N13468));
AOI22X1 inst_cellmath__50_0_I1289 (.Y(N5206), .A0(N5228), .A1(N5265), .B0(N5243), .B1(N5191));
AOI22X1 inst_cellmath__50_0_I8006 (.Y(N13523), .A0(N5135), .A1(N13540), .B0(N5206), .B1(N5171));
AOI22X1 inst_cellmath__50_0_I1290 (.Y(N5240), .A0(N5137), .A1(N5228), .B0(N5191), .B1(N5279));
AOI22X1 inst_cellmath__50_0_I8007 (.Y(inst_cellmath__50[10]), .A0(N5135), .A1(N13483), .B0(N5171), .B1(N5240));
AOI22X1 inst_cellmath__50_0_I8008 (.Y(inst_cellmath__50[11]), .A0(N13540), .A1(N5171), .B0(N13500), .B1(N5135));
AOI22X1 inst_cellmath__50_0_I8009 (.Y(inst_cellmath__50[12]), .A0(N5171), .A1(N13483), .B0(N5135), .B1(N13515));
OAI2BB1X1 inst_cellmath__50_0_I8154 (.Y(N13469), .A0N(N5228), .A1N(N13486), .B0(N13489));
INVX1 inst_cellmath__50_0_I8011 (.Y(N13485), .A(N13469));
AOI22X1 inst_cellmath__50_0_I8012 (.Y(N13512), .A0(N5135), .A1(N13485), .B0(N5171), .B1(N13500));
OAI2BB1X1 inst_cellmath__50_0_I8156 (.Y(N13513), .A0N(N5228), .A1N(N13504), .B0(N13499));
INVX1 inst_cellmath__50_0_I8014 (.Y(N13528), .A(N13513));
AOI22X1 inst_cellmath__50_0_I8015 (.Y(inst_cellmath__50[14]), .A0(N5135), .A1(N13528), .B0(N5171), .B1(N13515));
AOI22X1 inst_cellmath__50_0_I8016 (.Y(N13472), .A0(N5171), .A1(N13485), .B0(N5135), .B1(N5162));
AOI22X1 inst_cellmath__50_0_I8017 (.Y(inst_cellmath__50[16]), .A0(N5171), .A1(N13528), .B0(N5135), .B1(N5199));
INVXL buf1_A_I8290 (.Y(N13894), .A(N13523));
INVXL buf1_A_I8291 (.Y(inst_cellmath__50[9]), .A(N13894));
AND2XL inst_cellmath__50_0_I8019 (.Y(N5539), .A(inst_cellmath__50[10]), .B(inst_cellmath__50[9]));
INVXL buf1_A_I8292 (.Y(N13899), .A(N13512));
INVXL buf1_A_I8293 (.Y(inst_cellmath__50[13]), .A(N13899));
NAND2X1 inst_cellmath__50_0_I8023 (.Y(N13503), .A(N13523), .B(inst_cellmath__50[10]));
NOR2BX1 inst_cellmath__50_0_I8158 (.Y(N13479), .AN(inst_cellmath__50[12]), .B(N13503));
AND3XL inst_cellmath__50_0_I8025 (.Y(N5580), .A(inst_cellmath__50[11]), .B(inst_cellmath__50[12]), .C(N5539));
NAND2X1 inst_cellmath__50_0_I8026 (.Y(N13493), .A(N13472), .B(inst_cellmath__50[16]));
NAND2X1 inst_cellmath__50_0_I8027 (.Y(N13478), .A(N13512), .B(inst_cellmath__50[14]));
NAND2X1 inst_cellmath__50_0_I8028 (.Y(N13519), .A(inst_cellmath__50[11]), .B(N13479));
NOR3X2 inst_cellmath__50_0_I8029 (.Y(N5576), .A(N13493), .B(N13478), .C(N13519));
INVXL buf1_A_I8294 (.Y(N13904), .A(N13472));
INVXL buf1_A_I8295 (.Y(inst_cellmath__50[15]), .A(N13904));
MXI2XL inst_cellmath__50_0_I7869 (.Y(N13275), .A(N5139), .B(N13272), .S0(N5135));
AO22XL inst_cellmath__50_0_I7870 (.Y(inst_cellmath__50[2]), .A0(N5139), .A1(inst_cellmath__49[1]), .B0(N5135), .B1(N13272));
AOI22XL inst_cellmath__50_0_I7871 (.Y(inst_cellmath__50[3]), .A0(N5211), .A1(inst_cellmath__49[1]), .B0(N5189), .B1(N5135));
AOI22XL inst_cellmath__50_0_I7872 (.Y(inst_cellmath__50[4]), .A0(inst_cellmath__49[1]), .A1(N13272), .B0(N5135), .B1(N5261));
NOR2X1 inst_cellmath__50_0_I1310 (.Y(inst_cellmath__50[1]), .A(N5171), .B(N5211));
OR2XL cynw_cm_float_add2_ieee_I1337 (.Y(N628), .A(inst_cellmath__33[24]), .B(inst_cellmath__42));
XNOR2XL cynw_cm_float_add2_ieee_I1334 (.Y(N626), .A(inst_cellmath__42), .B(inst_cellmath__33[24]));
NOR2XL cynw_cm_float_add2_ieee_I1336 (.Y(N627), .A(N626), .B(inst_cellmath__30));
AO21XL cynw_cm_float_add2_ieee_I3005 (.Y(N630), .A0(inst_cellmath__30), .A1(N628), .B0(N627));
MX2XL cynw_cm_float_add2_ieee_I1340 (.Y(inst_cellmath__43), .A(inst_cellmath__33[24]), .B(N630), .S0(inst_cellmath__39[25]));
MXI2X1 inst_cellmath__50_0_I7873 (.Y(N13309), .A(inst_cellmath__50[1]), .B(inst_cellmath__43), .S0(inst_cellmath__49[1]));
NOR3BXL cynw_cm_float_add2_ieee_I1346 (.Y(inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3BXL cynw_cm_float_add2_ieee_I1342 (.Y(inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
NOR2BX1 cynw_cm_float_add2_ieee_I3006 (.Y(N635), .AN(inst_cellmath__5), .B(inst_cellmath__48));
AND2XL cynw_cm_float_add2_ieee_I1345 (.Y(N634), .A(inst_cellmath__6), .B(inst_cellmath__48));
NOR3XL cynw_cm_float_add2_ieee_I1347 (.Y(inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
OR2XL inst_cellmath__54__33__I1348 (.Y(N5486), .A(inst_cellmath__43), .B(inst_cellmath__42));
NOR2X2 inst_cellmath__50_0_I1309 (.Y(inst_cellmath__50[0]), .A(N5171), .B(N5139));
OR2XL inst_cellmath__54__33__I1349 (.Y(N631), .A(N5486), .B(inst_cellmath__50[0]));
MXI2XL cynw_cm_float_add2_ieee_I3104 (.Y(inst_cellmath__54), .A(N631), .B(inst_cellmath__42), .S0(inst_cellmath__49[1]));
NAND2XL cynw_cm_float_add2_ieee_I1351 (.Y(N632), .A(inst_cellmath__50[2]), .B(inst_cellmath__54));
CLKAND2X3 cynw_cm_float_add2_ieee_I1352 (.Y(N633), .A(inst_cellmath__4), .B(N632));
NOR4X2 inst_cellmath__50_0_I7874 (.Y(N13269), .A(N634), .B(N635), .C(inst_cellmath__8), .D(N633));
NOR2XL cynw_cm_float_add2_ieee_I1355 (.Y(N638), .A(N635), .B(N634));
NOR2XL inst_cellmath__50_0_I7875 (.Y(N13280), .A(N638), .B(inst_cellmath__54));
NOR2XL andori2bb1_A_I8296 (.Y(N13908), .A(N13309), .B(N13269));
NOR2XL andori2bb1_A_I8297 (.Y(inst_cellmath__55), .A(N13908), .B(N13280));
NOR2XL inst_cellmath__50_0_I7877 (.Y(N5600), .A(inst_cellmath__55), .B(inst_cellmath__50[2]));
NOR2X2 inst_cellmath__50_0_I7878 (.Y(N13312), .A(N13309), .B(N13269));
MXI2XL inst_cellmath__50_0_I7879 (.Y(N13268), .A(N13294), .B(N13298), .S0(inst_cellmath__49[1]));
INVXL inst_cellmath__50_0_I7880 (.Y(N13305), .A(inst_cellmath__50[4]));
OAI21X2 inst_cellmath__50_0_I7881 (.Y(N13314), .A0(N13280), .A1(N13312), .B0(N13275));
NOR3X4 inst_cellmath__50_0_I7882 (.Y(N5557), .A(N13268), .B(N13305), .C(N13314));
AOI22XL inst_cellmath__50_0_I1287 (.Y(N5132), .A0(N5228), .A1(N5193), .B0(N5174), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1288 (.Y(N5169), .A0(N5228), .A1(N5229), .B0(N5210), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1299 (.Y(N5233), .A0(N5228), .A1(N5129), .B0(N5274), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1300 (.Y(N5269), .A0(N5228), .A1(N5166), .B0(N5148), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1301 (.Y(N5141), .A0(N5228), .A1(N5204), .B0(N5181), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1302 (.Y(N5177), .A0(N5228), .A1(N5238), .B0(N5218), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1303 (.Y(N5213), .A0(N5228), .A1(N5274), .B0(N5253), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1304 (.Y(N5248), .A0(N5228), .A1(N5148), .B0(N5290), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1305 (.Y(N5284), .A0(N5228), .A1(N5181), .B0(N5161), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1306 (.Y(N5157), .A0(N5228), .A1(N5218), .B0(N5198), .B1(N5191));
AOI22XL inst_cellmath__50_0_I1314 (.Y(inst_cellmath__50[5]), .A0(N5135), .A1(N5132), .B0(N5189), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1315 (.Y(inst_cellmath__50[6]), .A0(N5135), .A1(N5169), .B0(N5261), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1316 (.Y(inst_cellmath__50[7]), .A0(N5135), .A1(N5206), .B0(N5132), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1317 (.Y(inst_cellmath__50[8]), .A0(N5135), .A1(N5240), .B0(N5169), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1326 (.Y(inst_cellmath__50[17]), .A0(N5135), .A1(N5233), .B0(N5162), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1327 (.Y(inst_cellmath__50[18]), .A0(N5135), .A1(N5269), .B0(N5199), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1328 (.Y(inst_cellmath__50[19]), .A0(N5135), .A1(N5141), .B0(N5233), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1329 (.Y(inst_cellmath__50[20]), .A0(N5135), .A1(N5177), .B0(N5269), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1330 (.Y(inst_cellmath__50[21]), .A0(N5135), .A1(N5213), .B0(N5141), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1331 (.Y(inst_cellmath__50[22]), .A0(N5135), .A1(N5248), .B0(N5177), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1332 (.Y(inst_cellmath__50[23]), .A0(N5135), .A1(N5284), .B0(N5213), .B1(N5171));
AOI22XL inst_cellmath__50_0_I1333 (.Y(inst_cellmath__50[24]), .A0(N5135), .A1(N5157), .B0(N5248), .B1(N5171));
AND2XL inst_cellmath__57_0_I1359 (.Y(N5546), .A(inst_cellmath__50[6]), .B(inst_cellmath__50[5]));
AND2XL inst_cellmath__57_0_I1362 (.Y(N5595), .A(inst_cellmath__50[18]), .B(inst_cellmath__50[17]));
NAND4X2 inst_cellmath__57_0_I2626 (.Y(N8072), .A(inst_cellmath__50[7]), .B(inst_cellmath__50[8]), .C(N5546), .D(N5557));
CLKINVX1 inst_cellmath__57_0_I2627 (.Y(N5588), .A(N8072));
CLKAND2X3 inst_cellmath__57_0_I1367 (.Y(N5596), .A(N5576), .B(N5588));
AND2XL inst_cellmath__57_0_I1368 (.Y(N5568), .A(N5580), .B(N5588));
NAND4X4 inst_cellmath__57_0_I2628 (.Y(N8080), .A(inst_cellmath__50[19]), .B(inst_cellmath__50[20]), .C(N5595), .D(N5596));
CLKINVX2 inst_cellmath__57_0_I2629 (.Y(N5543), .A(N8080));
AND2XL inst_cellmath__57_0_I1370 (.Y(N5594), .A(N5546), .B(N5557));
AND2XL inst_cellmath__57_0_I1371 (.Y(N5567), .A(N5539), .B(N5588));
AND3XL inst_cellmath__57_0_I8170 (.Y(N5542), .A(inst_cellmath__50[13]), .B(inst_cellmath__50[14]), .C(N5568));
AND2XL inst_cellmath__57_0_I1373 (.Y(N5591), .A(N5595), .B(N5596));
NAND3X2 inst_cellmath__57_0_I2630 (.Y(N8086), .A(inst_cellmath__50[21]), .B(inst_cellmath__50[22]), .C(N5543));
CLKINVX1 inst_cellmath__57_0_I2631 (.Y(N5564), .A(N8086));
NAND2XL inst_cellmath__57_0_I1375 (.Y(N5538), .A(inst_cellmath__50[3]), .B(N5600));
NAND2XL inst_cellmath__57_0_I1376 (.Y(N5587), .A(inst_cellmath__50[5]), .B(N5557));
NAND2XL inst_cellmath__57_0_I1377 (.Y(N5561), .A(inst_cellmath__50[7]), .B(N5594));
AND2XL inst_cellmath__57_0_I2632 (.Y(N8092), .A(inst_cellmath__50[9]), .B(N5588));
NAND2XL inst_cellmath__57_0_I1379 (.Y(N5583), .A(inst_cellmath__50[11]), .B(N5567));
NAND2XL inst_cellmath__57_0_I1380 (.Y(N5556), .A(inst_cellmath__50[13]), .B(N5568));
NAND2XL inst_cellmath__57_0_I1381 (.Y(N5532), .A(inst_cellmath__50[15]), .B(N5542));
NAND2XL inst_cellmath__57_0_I1382 (.Y(N5579), .A(inst_cellmath__50[17]), .B(N5596));
NAND2XL inst_cellmath__57_0_I1383 (.Y(N5553), .A(inst_cellmath__50[19]), .B(N5591));
AND2XL inst_cellmath__57_0_I2634 (.Y(N8098), .A(inst_cellmath__50[21]), .B(N5543));
NAND2XL inst_cellmath__57_0_I1385 (.Y(N5575), .A(inst_cellmath__50[23]), .B(N5564));
NAND3X2 inst_cellmath__57_0_I2647 (.Y(N8139), .A(inst_cellmath__50[23]), .B(inst_cellmath__50[24]), .C(N5564));
CLKINVX1 inst_cellmath__57_0_I2648 (.Y(inst_cellmath__57[23]), .A(N8139));
XOR2XL inst_cellmath__57_0_I1387 (.Y(inst_cellmath__57[0]), .A(inst_cellmath__50[2]), .B(inst_cellmath__55));
XOR2XL inst_cellmath__57_0_I1388 (.Y(inst_cellmath__57[1]), .A(N5600), .B(inst_cellmath__50[3]));
XNOR2X1 inst_cellmath__57_0_I1389 (.Y(inst_cellmath__57[2]), .A(N5538), .B(inst_cellmath__50[4]));
XOR2XL inst_cellmath__57_0_I1390 (.Y(inst_cellmath__57[3]), .A(N5557), .B(inst_cellmath__50[5]));
XNOR2X1 inst_cellmath__57_0_I1391 (.Y(inst_cellmath__57[4]), .A(N5587), .B(inst_cellmath__50[6]));
XOR2XL inst_cellmath__57_0_I1392 (.Y(inst_cellmath__57[5]), .A(N5594), .B(inst_cellmath__50[7]));
XNOR2X1 inst_cellmath__57_0_I1393 (.Y(inst_cellmath__57[6]), .A(N5561), .B(inst_cellmath__50[8]));
XOR2XL inst_cellmath__57_0_I3110 (.Y(inst_cellmath__57[7]), .A(N5588), .B(inst_cellmath__50[9]));
XOR2XL inst_cellmath__57_0_I3017 (.Y(inst_cellmath__57[8]), .A(N8092), .B(inst_cellmath__50[10]));
XOR2XL inst_cellmath__57_0_I1396 (.Y(inst_cellmath__57[9]), .A(N5567), .B(inst_cellmath__50[11]));
XNOR2X1 inst_cellmath__57_0_I1397 (.Y(inst_cellmath__57[10]), .A(N5583), .B(inst_cellmath__50[12]));
XOR2XL inst_cellmath__57_0_I1398 (.Y(inst_cellmath__57[11]), .A(N5568), .B(inst_cellmath__50[13]));
XNOR2X1 inst_cellmath__57_0_I1399 (.Y(inst_cellmath__57[12]), .A(N5556), .B(inst_cellmath__50[14]));
XOR2XL inst_cellmath__57_0_I1400 (.Y(inst_cellmath__57[13]), .A(N5542), .B(inst_cellmath__50[15]));
XNOR2X1 inst_cellmath__57_0_I1401 (.Y(inst_cellmath__57[14]), .A(N5532), .B(inst_cellmath__50[16]));
XOR2XL inst_cellmath__57_0_I1402 (.Y(inst_cellmath__57[15]), .A(N5596), .B(inst_cellmath__50[17]));
XNOR2X1 inst_cellmath__57_0_I1403 (.Y(inst_cellmath__57[16]), .A(N5579), .B(inst_cellmath__50[18]));
XOR2XL inst_cellmath__57_0_I1404 (.Y(inst_cellmath__57[17]), .A(N5591), .B(inst_cellmath__50[19]));
XNOR2X1 inst_cellmath__57_0_I1405 (.Y(inst_cellmath__57[18]), .A(N5553), .B(inst_cellmath__50[20]));
XOR2XL inst_cellmath__57_0_I3111 (.Y(inst_cellmath__57[19]), .A(N5543), .B(inst_cellmath__50[21]));
XOR2XL inst_cellmath__57_0_I3019 (.Y(inst_cellmath__57[20]), .A(N8098), .B(inst_cellmath__50[22]));
XOR2XL inst_cellmath__57_0_I3112 (.Y(inst_cellmath__57[21]), .A(N5564), .B(inst_cellmath__50[23]));
XNOR2X1 inst_cellmath__57_0_I1409 (.Y(inst_cellmath__57[22]), .A(N5575), .B(inst_cellmath__50[24]));
AO21XL cynw_cm_float_add2_ieee_I3113 (.Y(N642), .A0(inst_cellmath__45[24]), .A1(inst_cellmath__57[23]), .B0(inst_cellmath__45[25]));
INVXL buf1_A_I8298 (.Y(N13916), .A(N3367));
INVXL buf1_A_I8299 (.Y(N13433), .A(N13916));
INVXL inst_cellmath__59_0_I7919 (.Y(N574), .A(N13433));
MX2XL inst_cellmath__29_0_I1412 (.Y(inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(N574));
MX2XL inst_cellmath__29_0_I1413 (.Y(inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(N574));
MX2XL inst_cellmath__29_0_I1414 (.Y(inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(N574));
MX2XL inst_cellmath__29_0_I1415 (.Y(inst_cellmath__29[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(N574));
MX2XL inst_cellmath__29_0_I1416 (.Y(inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(N574));
MX2XL inst_cellmath__59_0_I7921 (.Y(inst_cellmath__29[6]), .A(b_exp[6]), .B(a_exp[6]), .S0(N13433));
MX2XL inst_cellmath__59_0_I7920 (.Y(inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(N574));
MX2XL inst_cellmath__59_0_I8080 (.Y(inst_cellmath__29[7]), .A(b_exp[7]), .B(a_exp[7]), .S0(N13433));
NAND3XL cynw_cm_float_add2_ieee_I1421 (.Y(N5708), .A(inst_cellmath__29[6]), .B(inst_cellmath__29[7]), .C(inst_cellmath__29[5]));
NOR2XL cynw_cm_float_add2_ieee_I1422 (.Y(N5707), .A(inst_cellmath__29[0]), .B(N5708));
INVXL inst_cellmath__59_0_I1431 (.Y(N5738), .A(inst_cellmath__29[1]));
ADDHX1 inst_cellmath__59_0_I1432 (.CO(N5743), .S(N5729), .A(inst_cellmath__29[1]), .B(inst_cellmath__29[2]));
ADDHX1 inst_cellmath__59_0_I1433 (.CO(N5716), .S(N5754), .A(inst_cellmath__29[3]), .B(N5743));
ADDHX1 inst_cellmath__59_0_I1434 (.CO(N5736), .S(N5724), .A(inst_cellmath__29[4]), .B(N5716));
INVXL inst_cellmath__59_0_I1435 (.Y(N5746), .A(inst_cellmath__29[5]));
INVXL inst_cellmath__59_0_I7923 (.Y(N13439), .A(inst_cellmath__29[6]));
INVXL inst_cellmath__59_0_I7924 (.Y(N13446), .A(inst_cellmath__29[7]));
NAND3XL inst_cellmath__59_0_I8074 (.Y(N13707), .A(inst_cellmath__29[4]), .B(inst_cellmath__29[3]), .C(N5707));
ADDFXL inst_cellmath__59_0_I8075 (.CO(N13744), .S(inst_cellmath__59[0]), .A(N5247), .B(inst_cellmath__29[0]), .CI(inst_cellmath__57[23]));
ADDFHXL inst_cellmath__59_0_I8076 (.CO(N13695), .S(inst_cellmath__59[1]), .A(N5135), .B(N5738), .CI(N13744));
ADDFHXL inst_cellmath__59_0_I8077 (.CO(N13732), .S(inst_cellmath__59[2]), .A(N5191), .B(N5729), .CI(N13695));
ADDFHXL inst_cellmath__59_0_I8078 (.CO(N13685), .S(inst_cellmath__59[3]), .A(N5754), .B(N5270), .CI(N13732));
ADDFHXL inst_cellmath__59_0_I8079 (.CO(N13722), .S(inst_cellmath__59[4]), .A(N5142), .B(N5724), .CI(N13685));
ADDFHXL inst_cellmath__59_0_I8081 (.CO(N13746), .S(inst_cellmath__59[5]), .A(N5736), .B(N5746), .CI(N13722));
ADDFHXL inst_cellmath__59_0_I8082 (.CO(N13697), .S(inst_cellmath__59[6]), .A(N13439), .B(inst_cellmath__29[5]), .CI(N13746));
ADDFHXL inst_cellmath__59_0_I8083 (.CO(N13734), .S(N13686), .A(inst_cellmath__29[6]), .B(N13446), .CI(N13697));
NOR2XL inst_cellmath__59_0_I8084 (.Y(N13740), .A(inst_cellmath__29[7]), .B(N13734));
INVX2 inst_cellmath__59_0_I8089 (.Y(N13699), .A(N13686));
OR4X1 inst_cellmath__59_0_I8090 (.Y(N13681), .A(N706), .B(inst_cellmath__17), .C(inst_cellmath__12), .D(inst_cellmath__63));
NAND3XL inst_cellmath__59_0_I8091 (.Y(N13754), .A(inst_cellmath__29[1]), .B(inst_cellmath__29[2]), .C(N642));
NOR2XL inst_cellmath__59_0_I8092 (.Y(inst_cellmath__62), .A(N13707), .B(N13754));
NOR4X4 inst_cellmath__59_0_I8093 (.Y(N13701), .A(N13681), .B(inst_cellmath__49[5]), .C(inst_cellmath__62), .D(N13740));
OR4X1 inst_cellmath__59_0_I8173 (.Y(N13719), .A(inst_cellmath__59[2]), .B(inst_cellmath__59[4]), .C(inst_cellmath__59[5]), .D(inst_cellmath__59[6]));
OR3XL inst_cellmath__59_0_I8219 (.Y(N13692), .A(inst_cellmath__59[0]), .B(inst_cellmath__59[1]), .C(inst_cellmath__59[3]));
INVXL inst_cellmath__59_0_I8096 (.Y(N13742), .A(inst_cellmath__29[7]));
INVX2 inst_cellmath__59_0_I8097 (.Y(N13710), .A(N13734));
NAND2X4 inst_cellmath__59_0_I8098 (.Y(N13730), .A(N13742), .B(N13710));
NOR2X1 inst_cellmath__59_0_I8099 (.Y(N13683), .A(N13742), .B(N13710));
INVX2 inst_cellmath__59_0_I8100 (.Y(N13738), .A(N13683));
NAND3X6 inst_cellmath__59_0_I8101 (.Y(N13706), .A(N13738), .B(N13730), .C(N13699));
OAI31X4 inst_cellmath__59_0_I8102 (.Y(inst_cellmath__71), .A0(N13719), .A1(N13692), .A2(N13706), .B0(N13701));
DLY1X1 inst_cellmath__59_0_I8103 (.Y(inst_cellmath__59[7]), .A(N13686));
OR4X1 cynw_cm_float_add2_ieee_I3024 (.Y(N650), .A(inst_cellmath__4), .B(inst_cellmath__8), .C(N635), .D(N634));
AND2XL cynw_cm_float_add2_ieee_I1460 (.Y(N651), .A(N650), .B(inst_cellmath__62));
OR4X1 cynw_cm_float_add2_ieee_I1461 (.Y(inst_cellmath__68[0]), .A(inst_cellmath__17), .B(inst_cellmath__12), .C(inst_cellmath__63), .D(N651));
OR4X1 inst_cellmath__72_0_I3025 (.Y(N5869), .A(inst_cellmath__12), .B(inst_cellmath__17), .C(inst_cellmath__63), .D(inst_cellmath__62));
CLKINVX4 inst_cellmath__72_0_I1465 (.Y(N5875), .A(inst_cellmath__71));
INVX1 inst_cellmath__72_0_I1466 (.Y(N5857), .A(N5875));
MX2XL inst_cellmath__72_0_I1467 (.Y(x[23]), .A(inst_cellmath__59[0]), .B(inst_cellmath__68[0]), .S0(N5857));
MX2XL inst_cellmath__72_0_I1468 (.Y(x[24]), .A(inst_cellmath__59[1]), .B(N5869), .S0(N5857));
MX2XL inst_cellmath__72_0_I1469 (.Y(x[25]), .A(inst_cellmath__59[2]), .B(N5869), .S0(N5857));
MX2XL inst_cellmath__72_0_I1470 (.Y(x[26]), .A(inst_cellmath__59[3]), .B(N5869), .S0(N5857));
MX2XL inst_cellmath__72_0_I1471 (.Y(x[27]), .A(inst_cellmath__59[4]), .B(N5869), .S0(N5857));
MX2XL inst_cellmath__72_0_I1472 (.Y(x[28]), .A(inst_cellmath__59[5]), .B(N5869), .S0(N5857));
MX2XL inst_cellmath__72_0_I1473 (.Y(x[29]), .A(inst_cellmath__59[6]), .B(N5869), .S0(N5857));
MX2XL inst_cellmath__72_0_I1474 (.Y(x[30]), .A(inst_cellmath__59[7]), .B(N5869), .S0(N5857));
NAND2XL inst_cellmath__7_0_I1475 (.Y(N5893), .A(rm[0]), .B(rm[1]));
NOR2XL inst_cellmath__7_0_I1476 (.Y(inst_cellmath__7), .A(rm[2]), .B(N5893));
XNOR2X1 cynw_cm_float_add2_ieee_I1477 (.Y(N652), .A(inst_cellmath__48), .B(inst_cellmath__5));
OR2XL cynw_cm_float_add2_ieee_I1478 (.Y(N653), .A(inst_cellmath__7), .B(N652));
NOR3BXL inst_cellmath__70_0_I1479 (.Y(N5912), .AN(N653), .B(inst_cellmath__8), .C(inst_cellmath__4));
AND2X1 inst_cellmath__70_0_I1480 (.Y(inst_cellmath__70), .A(inst_cellmath__62), .B(N5912));
CLKINVX4 inst_cellmath__73_0_I2919 (.Y(N8183), .A(N5875));
CLKINVX4 inst_cellmath__73_0_I2924 (.Y(N8188), .A(N8183));
INVXL inst_cellmath__73_0_I2922 (.Y(N8186), .A(N8183));
INVXL inst_cellmath__73_0_I2921 (.Y(N8185), .A(N8183));
INVXL inst_cellmath__73_0_I2920 (.Y(N8184), .A(N8183));
NOR2X6 inst_cellmath__73_0_I1482 (.Y(N5997), .A(inst_cellmath__63), .B(N5875));
NOR2BX4 inst_cellmath__73_0_I1483 (.Y(N5942), .AN(inst_cellmath__63), .B(N8188));
AOI22XL inst_cellmath__73_0_I1484 (.Y(N5926), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[0]));
AOI22XL inst_cellmath__73_0_I1485 (.Y(N5969), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[1]));
AOI22XL inst_cellmath__73_0_I1486 (.Y(N6011), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[2]));
AOI22XL inst_cellmath__73_0_I1487 (.Y(N5956), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[3]));
AOI22XL inst_cellmath__73_0_I1488 (.Y(N5999), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[4]));
AOI22XL inst_cellmath__73_0_I1489 (.Y(N5943), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[5]));
AOI22XL inst_cellmath__73_0_I1490 (.Y(N5986), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[6]));
AOI22XL inst_cellmath__73_0_I1491 (.Y(N5930), .A0(inst_cellmath__70), .A1(N5997), .B0(N8188), .B1(inst_cellmath__57[7]));
AOI22XL inst_cellmath__73_0_I1492 (.Y(N5973), .A0(inst_cellmath__70), .A1(N5997), .B0(N8186), .B1(inst_cellmath__57[8]));
AOI22XL inst_cellmath__73_0_I1493 (.Y(N5918), .A0(inst_cellmath__70), .A1(N5997), .B0(N8186), .B1(inst_cellmath__57[9]));
AOI22XL inst_cellmath__73_0_I1494 (.Y(N5961), .A0(inst_cellmath__70), .A1(N5997), .B0(N8186), .B1(inst_cellmath__57[10]));
AOI22XL inst_cellmath__73_0_I1495 (.Y(N6003), .A0(inst_cellmath__70), .A1(N5997), .B0(N8186), .B1(inst_cellmath__57[11]));
AOI22XL inst_cellmath__73_0_I1496 (.Y(N5947), .A0(inst_cellmath__70), .A1(N5997), .B0(N8186), .B1(inst_cellmath__57[12]));
AOI22XL inst_cellmath__73_0_I1497 (.Y(N5990), .A0(inst_cellmath__70), .A1(N5997), .B0(N8185), .B1(inst_cellmath__57[13]));
AOI22XL inst_cellmath__73_0_I1498 (.Y(N5934), .A0(inst_cellmath__70), .A1(N5997), .B0(N8185), .B1(inst_cellmath__57[14]));
AOI22XL inst_cellmath__73_0_I1499 (.Y(N5978), .A0(inst_cellmath__70), .A1(N5997), .B0(N8185), .B1(inst_cellmath__57[15]));
AOI22XL inst_cellmath__73_0_I1500 (.Y(N5923), .A0(inst_cellmath__70), .A1(N5997), .B0(N8185), .B1(inst_cellmath__57[16]));
AOI22XL inst_cellmath__73_0_I1501 (.Y(N5966), .A0(inst_cellmath__70), .A1(N5997), .B0(N8185), .B1(inst_cellmath__57[17]));
AOI22XL inst_cellmath__73_0_I1502 (.Y(N6008), .A0(inst_cellmath__70), .A1(N5997), .B0(N8184), .B1(inst_cellmath__57[18]));
AOI22XL inst_cellmath__73_0_I1503 (.Y(N5953), .A0(inst_cellmath__70), .A1(N5997), .B0(N8184), .B1(inst_cellmath__57[19]));
AOI22XL inst_cellmath__73_0_I1504 (.Y(N5995), .A0(inst_cellmath__70), .A1(N5997), .B0(N8184), .B1(inst_cellmath__57[20]));
AOI22XL inst_cellmath__73_0_I1505 (.Y(N5939), .A0(inst_cellmath__70), .A1(N5997), .B0(N8184), .B1(inst_cellmath__57[21]));
AOI22XL inst_cellmath__73_0_I1506 (.Y(N5982), .A0(inst_cellmath__70), .A1(N5997), .B0(N8184), .B1(inst_cellmath__57[22]));
OAI2BB1XL inst_cellmath__73_0_I1507 (.Y(x[0]), .A0N(N5942), .A1N(inst_cellmath__64[0]), .B0(N5926));
OAI2BB1XL inst_cellmath__73_0_I1508 (.Y(x[1]), .A0N(N5942), .A1N(inst_cellmath__64[1]), .B0(N5969));
OAI2BB1XL inst_cellmath__73_0_I1509 (.Y(x[2]), .A0N(N5942), .A1N(inst_cellmath__64[2]), .B0(N6011));
OAI2BB1XL inst_cellmath__73_0_I1510 (.Y(x[3]), .A0N(N5942), .A1N(inst_cellmath__64[3]), .B0(N5956));
OAI2BB1XL inst_cellmath__73_0_I1511 (.Y(x[4]), .A0N(N5942), .A1N(inst_cellmath__64[4]), .B0(N5999));
OAI2BB1XL inst_cellmath__73_0_I1512 (.Y(x[5]), .A0N(N5942), .A1N(inst_cellmath__64[5]), .B0(N5943));
OAI2BB1XL inst_cellmath__73_0_I1513 (.Y(x[6]), .A0N(N5942), .A1N(inst_cellmath__64[6]), .B0(N5986));
OAI2BB1XL inst_cellmath__73_0_I1514 (.Y(x[7]), .A0N(N5942), .A1N(inst_cellmath__64[7]), .B0(N5930));
OAI2BB1XL inst_cellmath__73_0_I1515 (.Y(x[8]), .A0N(N5942), .A1N(inst_cellmath__64[8]), .B0(N5973));
OAI2BB1XL inst_cellmath__73_0_I1516 (.Y(x[9]), .A0N(N5942), .A1N(inst_cellmath__64[9]), .B0(N5918));
OAI2BB1XL inst_cellmath__73_0_I1517 (.Y(x[10]), .A0N(N5942), .A1N(inst_cellmath__64[10]), .B0(N5961));
OAI2BB1XL inst_cellmath__73_0_I1518 (.Y(x[11]), .A0N(N5942), .A1N(inst_cellmath__64[11]), .B0(N6003));
OAI2BB1XL inst_cellmath__73_0_I1519 (.Y(x[12]), .A0N(N5942), .A1N(inst_cellmath__64[12]), .B0(N5947));
OAI2BB1XL inst_cellmath__73_0_I1520 (.Y(x[13]), .A0N(N5942), .A1N(inst_cellmath__64[13]), .B0(N5990));
OAI2BB1XL inst_cellmath__73_0_I1521 (.Y(x[14]), .A0N(N5942), .A1N(inst_cellmath__64[14]), .B0(N5934));
OAI2BB1XL inst_cellmath__73_0_I1522 (.Y(x[15]), .A0N(N5942), .A1N(inst_cellmath__64[15]), .B0(N5978));
OAI2BB1XL inst_cellmath__73_0_I1523 (.Y(x[16]), .A0N(N5942), .A1N(inst_cellmath__64[16]), .B0(N5923));
OAI2BB1XL inst_cellmath__73_0_I1524 (.Y(x[17]), .A0N(N5942), .A1N(inst_cellmath__64[17]), .B0(N5966));
OAI2BB1XL inst_cellmath__73_0_I1525 (.Y(x[18]), .A0N(N5942), .A1N(inst_cellmath__64[18]), .B0(N6008));
OAI2BB1XL inst_cellmath__73_0_I1526 (.Y(x[19]), .A0N(N5942), .A1N(inst_cellmath__64[19]), .B0(N5953));
OAI2BB1XL inst_cellmath__73_0_I1527 (.Y(x[20]), .A0N(N5942), .A1N(inst_cellmath__64[20]), .B0(N5995));
OAI2BB1XL inst_cellmath__73_0_I1528 (.Y(x[21]), .A0N(N5942), .A1N(inst_cellmath__64[21]), .B0(N5939));
NAND2BXL inst_cellmath__73_0_I1529 (.Y(x[22]), .AN(N5942), .B(N5982));
assign inst_cellmath__27[0] = 1'B0;
assign inst_cellmath__33[0] = 1'B0;
assign inst_cellmath__33[1] = 1'B0;
assign inst_cellmath__33[2] = 1'B0;
assign inst_cellmath__33[3] = 1'B0;
assign inst_cellmath__33[4] = 1'B0;
assign inst_cellmath__33[5] = 1'B0;
assign inst_cellmath__33[6] = 1'B0;
assign inst_cellmath__33[7] = 1'B0;
assign inst_cellmath__33[8] = 1'B0;
assign inst_cellmath__33[9] = 1'B0;
assign inst_cellmath__33[10] = 1'B0;
assign inst_cellmath__33[11] = 1'B0;
assign inst_cellmath__33[12] = 1'B0;
assign inst_cellmath__33[13] = 1'B0;
assign inst_cellmath__33[14] = 1'B0;
assign inst_cellmath__33[15] = 1'B0;
assign inst_cellmath__33[16] = 1'B0;
assign inst_cellmath__33[17] = 1'B0;
assign inst_cellmath__33[18] = 1'B0;
assign inst_cellmath__33[19] = 1'B0;
assign inst_cellmath__33[20] = 1'B0;
assign inst_cellmath__33[21] = 1'B0;
assign inst_cellmath__33[22] = 1'B0;
assign inst_cellmath__33[23] = 1'B0;
assign inst_cellmath__33[27] = 1'B0;
assign inst_cellmath__33[28] = 1'B0;
assign inst_cellmath__33[31] = 1'B0;
assign inst_cellmath__33[32] = 1'B0;
assign inst_cellmath__33[33] = 1'B0;
assign inst_cellmath__33[36] = 1'B0;
assign inst_cellmath__33[37] = 1'B0;
assign inst_cellmath__33[41] = 1'B0;
assign inst_cellmath__36[0] = 1'B0;
assign inst_cellmath__36[1] = 1'B0;
assign inst_cellmath__36[2] = 1'B0;
assign inst_cellmath__36[3] = 1'B0;
assign inst_cellmath__36[4] = 1'B0;
assign inst_cellmath__36[5] = 1'B0;
assign inst_cellmath__36[6] = 1'B0;
assign inst_cellmath__36[7] = 1'B0;
assign inst_cellmath__36[8] = 1'B0;
assign inst_cellmath__36[9] = 1'B0;
assign inst_cellmath__36[10] = 1'B0;
assign inst_cellmath__36[11] = 1'B0;
assign inst_cellmath__36[12] = 1'B0;
assign inst_cellmath__36[13] = 1'B0;
assign inst_cellmath__36[14] = 1'B0;
assign inst_cellmath__36[15] = 1'B0;
assign inst_cellmath__36[16] = 1'B0;
assign inst_cellmath__36[17] = 1'B0;
assign inst_cellmath__36[18] = 1'B0;
assign inst_cellmath__36[19] = 1'B0;
assign inst_cellmath__36[20] = 1'B0;
assign inst_cellmath__36[21] = 1'B0;
assign inst_cellmath__36[22] = 1'B0;
assign inst_cellmath__36[23] = 1'B0;
assign inst_cellmath__36[24] = 1'B0;
assign inst_cellmath__36[25] = 1'B0;
assign inst_cellmath__36[49] = 1'B1;
assign inst_cellmath__37[1] = 1'B0;
assign inst_cellmath__37[2] = 1'B0;
assign inst_cellmath__37[42] = 1'B0;
assign inst_cellmath__37[45] = 1'B0;
assign inst_cellmath__37[46] = 1'B0;
assign inst_cellmath__37[47] = 1'B0;
assign inst_cellmath__37[48] = 1'B0;
assign inst_cellmath__37[49] = 1'B0;
assign inst_cellmath__39[2] = 1'B0;
assign inst_cellmath__39[3] = 1'B0;
assign inst_cellmath__39[5] = 1'B0;
assign inst_cellmath__39[6] = 1'B0;
assign inst_cellmath__39[24] = 1'B0;
assign inst_cellmath__45[26] = 1'B0;
assign inst_cellmath__49[2] = 1'B0;
assign inst_cellmath__49[3] = 1'B0;
assign inst_cellmath__49[4] = 1'B0;
assign inst_cellmath__59[8] = 1'B0;
assign inst_cellmath__59[9] = 1'B0;
assign inst_cellmath__64[22] = 1'B1;
assign inst_cellmath__68[1] = 1'B0;
assign inst_cellmath__68[2] = 1'B0;
assign inst_cellmath__68[3] = 1'B0;
assign inst_cellmath__68[4] = 1'B0;
assign inst_cellmath__68[5] = 1'B0;
assign inst_cellmath__68[6] = 1'B0;
assign inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  urL3TgrXqhA= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



