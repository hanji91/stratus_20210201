/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:38:04 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_5_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__71,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4838,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4917,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13685,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13732,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13740,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916;
wire N5507,N5514,N5521,N5528,N5535,N5542,N5549 
	,N5556,N5563,N5570,N5577,N5584,N5591,N5598,N5605 
	,N5612,N5619,N5626,N5633,N5640,N5647,N5654,N5718 
	,N5720,N5956,N5972,N5974,N5998,N6000,N6007,N6014 
	,N6021,N6028,N6035,N6042,N6049,N6056,N6063,N6070 
	,N6077,N6084,N6091,N6098,N6105,N6112,N6119,N6126 
	,N6133,N6140,N6147,N6154,N6299,N6304,N6430,N6439 
	,N6448,N6457,N6466,N6475,N6484,N6493,N6502,N6511 
	,N6520,N6529,N6538,N6547,N6565,N6574,N6583,N6592 
	,N6601,N6655,N6671,N6673,N6837,N6842,N6946,N7014 
	,N7038,N7040,N7068,N7070,N7083,N7091,N7099,N7128 
	,N7139,N7141,N7149,N7151,N7158,N7167,N7169,N7185 
	,N7187,N7203,N7205,N7221,N7223,N7230,N7239,N7241 
	,N7248,N7257,N7259,N7270,N7272,N7427,N7429,N7501 
	,N7505,N7661,N7663,N7931,N7933,N8017,N8100,N8102 
	,N8104,N8110,N8203,N8480,N8521,N8528,N8536,N8578 
	,N8941,N8990,N9246,N9251,N9260,N9267,N9274,N9281 
	,N9288,N9295,N9302,N9310,N9318,N9326,N9334,N9342 
	,N9350,N9358,N9366,N9374,N9382,N9390,N9398,N9404 
	,N9406,N9422,N9431,N9433,N9437,N9445,N9453,N9461 
	,N9469,N9477,N9485,N9493,N9501,N9509,N9517,N9525 
	,N9533,N9541,N9549,N9557,N9565,N9576,N10111,N10116 
	,N10123,N10157,N10159,N10166,N10168,N10173,N10175,N10193 
	,N10610,N10611,N10666,N10671;
reg x_reg_L1_12__retimed_I5171_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5171_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23];
	end
assign N10193 = x_reg_L1_12__retimed_I5171_QOUT;
reg x_reg_L1_14__retimed_I5162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5162_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14];
	end
assign N10175 = x_reg_L1_14__retimed_I5162_QOUT;
reg x_reg_L1_20__retimed_I5161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5161_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20];
	end
assign N10173 = x_reg_L1_20__retimed_I5161_QOUT;
reg x_reg_L0_22__retimed_I5159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5159_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627;
	end
assign N10168 = x_reg_L0_22__retimed_I5159_QOUT;
reg x_reg_L0_22__retimed_I5158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5158_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596;
	end
assign N10166 = x_reg_L0_22__retimed_I5158_QOUT;
reg x_reg_L0_22__retimed_I5156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5156_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684;
	end
assign N10159 = x_reg_L0_22__retimed_I5156_QOUT;
reg x_reg_L0_22__retimed_I5155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5155_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706;
	end
assign N10157 = x_reg_L0_22__retimed_I5155_QOUT;
reg x_reg_L0_22__retimed_I5141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5141_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3];
	end
assign N10123 = x_reg_L0_22__retimed_I5141_QOUT;
reg x_reg_L0_22__retimed_I5139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5139_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7];
	end
assign N10116 = x_reg_L0_22__retimed_I5139_QOUT;
reg x_reg_L0_22__retimed_I5137_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5137_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4];
	end
assign N10111 = x_reg_L0_22__retimed_I5137_QOUT;
reg x_reg_L0_22__retimed_I4892_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4892_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621;
	end
assign N9576 = x_reg_L0_22__retimed_I4892_QOUT;
reg x_reg_L0_22__retimed_I4888_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4888_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719;
	end
assign N9565 = x_reg_L0_22__retimed_I4888_QOUT;
reg x_reg_L0_22__retimed_I4885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4885_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647;
	end
assign N9557 = x_reg_L0_22__retimed_I4885_QOUT;
reg x_reg_L0_22__retimed_I4882_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4882_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579;
	end
assign N9549 = x_reg_L0_22__retimed_I4882_QOUT;
reg x_reg_L0_22__retimed_I4879_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4879_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653;
	end
assign N9541 = x_reg_L0_22__retimed_I4879_QOUT;
reg x_reg_L0_22__retimed_I4876_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4876_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589;
	end
assign N9533 = x_reg_L0_22__retimed_I4876_QOUT;
reg x_reg_L0_22__retimed_I4873_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4873_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663;
	end
assign N9525 = x_reg_L0_22__retimed_I4873_QOUT;
reg x_reg_L0_22__retimed_I4870_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4870_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595;
	end
assign N9517 = x_reg_L0_22__retimed_I4870_QOUT;
reg x_reg_L0_22__retimed_I4867_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4867_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673;
	end
assign N9509 = x_reg_L0_22__retimed_I4867_QOUT;
reg x_reg_L0_22__retimed_I4864_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4864_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603;
	end
assign N9501 = x_reg_L0_22__retimed_I4864_QOUT;
reg x_reg_L0_22__retimed_I4861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4861_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679;
	end
assign N9493 = x_reg_L0_22__retimed_I4861_QOUT;
reg x_reg_L0_22__retimed_I4858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4858_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609;
	end
assign N9485 = x_reg_L0_22__retimed_I4858_QOUT;
reg x_reg_L0_22__retimed_I4855_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4855_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687;
	end
assign N9477 = x_reg_L0_22__retimed_I4855_QOUT;
reg x_reg_L0_22__retimed_I4852_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4852_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618;
	end
assign N9469 = x_reg_L0_22__retimed_I4852_QOUT;
reg x_reg_L0_22__retimed_I4849_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4849_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695;
	end
assign N9461 = x_reg_L0_22__retimed_I4849_QOUT;
reg x_reg_L0_22__retimed_I4846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4846_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626;
	end
assign N9453 = x_reg_L0_22__retimed_I4846_QOUT;
reg x_reg_L0_22__retimed_I4843_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4843_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704;
	end
assign N9445 = x_reg_L0_22__retimed_I4843_QOUT;
reg x_reg_L0_22__retimed_I4840_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4840_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257;
	end
assign N9437 = x_reg_L0_22__retimed_I4840_QOUT;
reg x_reg_L0_22__retimed_I4839_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4839_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634;
	end
assign N9433 = x_reg_L0_22__retimed_I4839_QOUT;
reg x_reg_L0_22__retimed_I4838_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4838_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613;
	end
assign N9431 = x_reg_L0_22__retimed_I4838_QOUT;
reg x_reg_L0_22__retimed_I4834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4834_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604;
	end
assign N9422 = x_reg_L0_22__retimed_I4834_QOUT;
reg x_reg_L0_22__retimed_I4829_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4829_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604;
	end
assign N9406 = x_reg_L0_22__retimed_I4829_QOUT;
reg x_reg_L0_22__retimed_I4828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4828_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667;
	end
assign N9404 = x_reg_L0_22__retimed_I4828_QOUT;
reg x_reg_L0_22__retimed_I4827_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4827_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586;
	end
assign N9398 = x_reg_L0_22__retimed_I4827_QOUT;
reg x_reg_L0_22__retimed_I4825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4825_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668;
	end
assign N9390 = x_reg_L0_22__retimed_I4825_QOUT;
reg x_reg_L0_22__retimed_I4823_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4823_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648;
	end
assign N9382 = x_reg_L0_22__retimed_I4823_QOUT;
reg x_reg_L0_22__retimed_I4821_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4821_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713;
	end
assign N9374 = x_reg_L0_22__retimed_I4821_QOUT;
reg x_reg_L0_22__retimed_I4819_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4819_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628;
	end
assign N9366 = x_reg_L0_22__retimed_I4819_QOUT;
reg x_reg_L0_22__retimed_I4817_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4817_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692;
	end
assign N9358 = x_reg_L0_22__retimed_I4817_QOUT;
reg x_reg_L0_22__retimed_I4815_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4815_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610;
	end
assign N9350 = x_reg_L0_22__retimed_I4815_QOUT;
reg x_reg_L0_22__retimed_I4813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4813_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676;
	end
assign N9342 = x_reg_L0_22__retimed_I4813_QOUT;
reg x_reg_L0_22__retimed_I4811_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4811_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593;
	end
assign N9334 = x_reg_L0_22__retimed_I4811_QOUT;
reg x_reg_L0_22__retimed_I4809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4809_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654;
	end
assign N9326 = x_reg_L0_22__retimed_I4809_QOUT;
reg x_reg_L0_22__retimed_I4807_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4807_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722;
	end
assign N9318 = x_reg_L0_22__retimed_I4807_QOUT;
reg x_reg_L0_22__retimed_I4805_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4805_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636;
	end
assign N9310 = x_reg_L0_22__retimed_I4805_QOUT;
reg x_reg_L0_22__retimed_I4803_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4803_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700;
	end
assign N9302 = x_reg_L0_22__retimed_I4803_QOUT;
reg x_reg_L0_22__retimed_I4801_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4801_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620;
	end
assign N9295 = x_reg_L0_22__retimed_I4801_QOUT;
reg x_reg_L0_22__retimed_I4799_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4799_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682;
	end
assign N9288 = x_reg_L0_22__retimed_I4799_QOUT;
reg x_reg_L0_22__retimed_I4797_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4797_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600;
	end
assign N9281 = x_reg_L0_22__retimed_I4797_QOUT;
reg x_reg_L0_22__retimed_I4795_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4795_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665;
	end
assign N9274 = x_reg_L0_22__retimed_I4795_QOUT;
reg x_reg_L0_22__retimed_I4793_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4793_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582;
	end
assign N9267 = x_reg_L0_22__retimed_I4793_QOUT;
reg x_reg_L0_22__retimed_I4791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4791_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644;
	end
assign N9260 = x_reg_L0_22__retimed_I4791_QOUT;
reg x_reg_L0_22__retimed_I4788_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4788_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
	end
assign N9251 = x_reg_L0_22__retimed_I4788_QOUT;
reg x_reg_L0_22__retimed_I4787_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4787_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677;
	end
assign N9246 = x_reg_L0_22__retimed_I4787_QOUT;
reg x_reg_L0_22__retimed_I4696_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4696_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848;
	end
assign N8990 = x_reg_L0_22__retimed_I4696_QOUT;
reg x_reg_L0_22__retimed_I4678_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4678_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827;
	end
assign N8941 = x_reg_L0_22__retimed_I4678_QOUT;
reg x_reg_L0_22__retimed_I4607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4607_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486;
	end
assign N8578 = x_reg_L0_22__retimed_I4607_QOUT;
reg x_reg_L0_22__retimed_I4593_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4593_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N8536 = x_reg_L0_22__retimed_I4593_QOUT;
reg x_reg_L0_22__retimed_I4590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4590_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N8528 = x_reg_L0_22__retimed_I4590_QOUT;
reg x_reg_L0_22__retimed_I4587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4587_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N8521 = x_reg_L0_22__retimed_I4587_QOUT;
reg x_reg_L0_22__retimed_I4570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4570_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
	end
assign N8480 = x_reg_L0_22__retimed_I4570_QOUT;
reg x_reg_L0_22__retimed_I4480_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4480_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4;
	end
assign N8203 = x_reg_L0_22__retimed_I4480_QOUT;
reg x_reg_L0_22__retimed_I4443_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4443_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43;
	end
assign N8110 = x_reg_L0_22__retimed_I4443_QOUT;
reg x_reg_L0_22__retimed_I4441_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4441_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N8104 = x_reg_L0_22__retimed_I4441_QOUT;
reg x_reg_L0_22__retimed_I4440_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4440_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635;
	end
assign N8102 = x_reg_L0_22__retimed_I4440_QOUT;
reg x_reg_L0_22__retimed_I4439_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4439_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
	end
assign N8100 = x_reg_L0_22__retimed_I4439_QOUT;
reg x_reg_L0_22__retimed_I4406_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4406_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638;
	end
assign N8017 = x_reg_L0_22__retimed_I4406_QOUT;
reg x_reg_L1_21__retimed_I4373_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I4373_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23];
	end
assign N7933 = x_reg_L1_21__retimed_I4373_QOUT;
reg x_reg_L1_21__retimed_I4372_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I4372_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564;
	end
assign N7931 = x_reg_L1_21__retimed_I4372_QOUT;
reg x_reg_L1_22__retimed_I4270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I4270_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24];
	end
assign N7663 = x_reg_L1_22__retimed_I4270_QOUT;
reg x_reg_L1_22__retimed_I4269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I4269_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575;
	end
assign N7661 = x_reg_L1_22__retimed_I4269_QOUT;
reg x_reg_L1_12__retimed_I4208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4208_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
	end
assign N7505 = x_reg_L1_12__retimed_I4208_QOUT;
reg x_reg_L1_12__retimed_I4206_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4206_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24];
	end
assign N7501 = x_reg_L1_12__retimed_I4206_QOUT;
reg x_reg_L1_12__retimed_I4178_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4178_QOUT <= N7070;
	end
assign N7429 = x_reg_L1_12__retimed_I4178_QOUT;
reg x_reg_L1_12__retimed_I4177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4177_QOUT <= N7068;
	end
assign N7427 = x_reg_L1_12__retimed_I4177_QOUT;
reg x_reg_L1_23__retimed_I4115_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I4115_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247;
	end
assign N7272 = x_reg_L1_23__retimed_I4115_QOUT;
reg x_reg_L1_23__retimed_I4114_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I4114_QOUT <= N7248;
	end
assign N7270 = x_reg_L1_23__retimed_I4114_QOUT;
reg x_reg_L1_24__retimed_I4111_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I4111_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135;
	end
assign N7259 = x_reg_L1_24__retimed_I4111_QOUT;
reg x_reg_L1_24__retimed_I4110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I4110_QOUT <= N7230;
	end
assign N7257 = x_reg_L1_24__retimed_I4110_QOUT;
reg x_reg_L0_22__retimed_I4107_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4107_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0];
	end
assign N7248 = x_reg_L0_22__retimed_I4107_QOUT;
reg x_reg_L1_25__retimed_I4105_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I4105_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191;
	end
assign N7241 = x_reg_L1_25__retimed_I4105_QOUT;
reg x_reg_L1_25__retimed_I4104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I4104_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729;
	end
assign N7239 = x_reg_L1_25__retimed_I4104_QOUT;
reg x_reg_L0_22__retimed_I4101_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4101_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738;
	end
assign N7230 = x_reg_L0_22__retimed_I4101_QOUT;
reg x_reg_L1_26__retimed_I4099_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I4099_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754;
	end
assign N7223 = x_reg_L1_26__retimed_I4099_QOUT;
reg x_reg_L1_26__retimed_I4098_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I4098_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270;
	end
assign N7221 = x_reg_L1_26__retimed_I4098_QOUT;
reg x_reg_L1_27__retimed_I4093_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I4093_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142;
	end
assign N7205 = x_reg_L1_27__retimed_I4093_QOUT;
reg x_reg_L1_27__retimed_I4092_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I4092_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724;
	end
assign N7203 = x_reg_L1_27__retimed_I4092_QOUT;
reg x_reg_L1_28__retimed_I4087_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I4087_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736;
	end
assign N7187 = x_reg_L1_28__retimed_I4087_QOUT;
reg x_reg_L1_28__retimed_I4086_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I4086_QOUT <= N7158;
	end
assign N7185 = x_reg_L1_28__retimed_I4086_QOUT;
reg x_reg_L1_29__retimed_I4081_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I4081_QOUT <= N7141;
	end
assign N7169 = x_reg_L1_29__retimed_I4081_QOUT;
reg x_reg_L1_29__retimed_I4080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I4080_QOUT <= N7139;
	end
assign N7167 = x_reg_L1_29__retimed_I4080_QOUT;
reg x_reg_L0_22__retimed_I4077_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4077_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
	end
assign N7158 = x_reg_L0_22__retimed_I4077_QOUT;
reg x_reg_L1_30__retimed_I4075_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I4075_QOUT <= N7128;
	end
assign N7151 = x_reg_L1_30__retimed_I4075_QOUT;
reg x_reg_L1_30__retimed_I4074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I4074_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446;
	end
assign N7149 = x_reg_L1_30__retimed_I4074_QOUT;
reg x_reg_L0_22__retimed_I4072_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4072_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439;
	end
assign N7141 = x_reg_L0_22__retimed_I4072_QOUT;
reg x_reg_L0_22__retimed_I4071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4071_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
	end
assign N7139 = x_reg_L0_22__retimed_I4071_QOUT;
reg x_reg_L0_22__retimed_I4068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4068_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
	end
assign N7128 = x_reg_L0_22__retimed_I4068_QOUT;
reg x_reg_L1_12__retimed_I4058_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4058_QOUT <= N7014;
	end
assign N7099 = x_reg_L1_12__retimed_I4058_QOUT;
reg x_reg_L1_12__retimed_I4056_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4056_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742;
	end
assign N7091 = x_reg_L1_12__retimed_I4056_QOUT;
reg x_reg_L1_12__retimed_I4053_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4053_QOUT <= N10116;
	end
assign N7083 = x_reg_L1_12__retimed_I4053_QOUT;
reg x_reg_L0_22__retimed_I4049_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4049_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2];
	end
assign N7070 = x_reg_L0_22__retimed_I4049_QOUT;
reg x_reg_L0_22__retimed_I4048_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4048_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
	end
assign N7068 = x_reg_L0_22__retimed_I4048_QOUT;
reg x_reg_L1_12__retimed_I4036_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4036_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5];
	end
assign N7040 = x_reg_L1_12__retimed_I4036_QOUT;
reg x_reg_L1_12__retimed_I4035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4035_QOUT <= N6946;
	end
assign N7038 = x_reg_L1_12__retimed_I4035_QOUT;
reg x_reg_L0_22__retimed_I4026_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4026_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707;
	end
assign N7014 = x_reg_L0_22__retimed_I4026_QOUT;
reg x_reg_L0_22__retimed_I3999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3999_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681;
	end
assign N6946 = x_reg_L0_22__retimed_I3999_QOUT;
reg x_reg_L1_23__retimed_I3965_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3965_QOUT <= N6304;
	end
assign N6842 = x_reg_L1_23__retimed_I3965_QOUT;
reg x_reg_L1_22__retimed_I3963_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I3963_QOUT <= N6299;
	end
assign N6837 = x_reg_L1_22__retimed_I3963_QOUT;
reg x_reg_L1_23__retimed_I3927_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3927_QOUT <= N5974;
	end
assign N6673 = x_reg_L1_23__retimed_I3927_QOUT;
reg x_reg_L1_23__retimed_I3926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3926_QOUT <= N5972;
	end
assign N6671 = x_reg_L1_23__retimed_I3926_QOUT;
reg x_reg_L1_22__retimed_I3923_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I3923_QOUT <= N5956;
	end
assign N6655 = x_reg_L1_22__retimed_I3923_QOUT;
reg x_reg_L1_19__retimed_I3909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3909_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19];
	end
assign N6601 = x_reg_L1_19__retimed_I3909_QOUT;
reg x_reg_L1_18__retimed_I3905_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3905_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18];
	end
assign N6592 = x_reg_L1_18__retimed_I3905_QOUT;
reg x_reg_L1_17__retimed_I3901_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3901_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17];
	end
assign N6583 = x_reg_L1_17__retimed_I3901_QOUT;
reg x_reg_L1_16__retimed_I3897_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3897_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16];
	end
assign N6574 = x_reg_L1_16__retimed_I3897_QOUT;
reg x_reg_L1_15__retimed_I3893_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3893_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15];
	end
assign N6565 = x_reg_L1_15__retimed_I3893_QOUT;
reg x_reg_L1_13__retimed_I3885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3885_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13];
	end
assign N6547 = x_reg_L1_13__retimed_I3885_QOUT;
reg x_reg_L1_12__retimed_I3881_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3881_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12];
	end
assign N6538 = x_reg_L1_12__retimed_I3881_QOUT;
reg x_reg_L1_11__retimed_I3877_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I3877_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11];
	end
assign N6529 = x_reg_L1_11__retimed_I3877_QOUT;
reg x_reg_L1_10__retimed_I3873_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I3873_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10];
	end
assign N6520 = x_reg_L1_10__retimed_I3873_QOUT;
reg x_reg_L1_9__retimed_I3869_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I3869_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9];
	end
assign N6511 = x_reg_L1_9__retimed_I3869_QOUT;
reg x_reg_L1_8__retimed_I3865_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3865_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8];
	end
assign N6502 = x_reg_L1_8__retimed_I3865_QOUT;
reg x_reg_L1_7__retimed_I3861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3861_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7];
	end
assign N6493 = x_reg_L1_7__retimed_I3861_QOUT;
reg x_reg_L1_6__retimed_I3857_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3857_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6];
	end
assign N6484 = x_reg_L1_6__retimed_I3857_QOUT;
reg x_reg_L1_5__retimed_I3853_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3853_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5];
	end
assign N6475 = x_reg_L1_5__retimed_I3853_QOUT;
reg x_reg_L1_4__retimed_I3849_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3849_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4];
	end
assign N6466 = x_reg_L1_4__retimed_I3849_QOUT;
reg x_reg_L1_3__retimed_I3845_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3845_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3];
	end
assign N6457 = x_reg_L1_3__retimed_I3845_QOUT;
reg x_reg_L1_2__retimed_I3841_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3841_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2];
	end
assign N6448 = x_reg_L1_2__retimed_I3841_QOUT;
reg x_reg_L1_1__retimed_I3837_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3837_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1];
	end
assign N6439 = x_reg_L1_1__retimed_I3837_QOUT;
reg x_reg_L1_0__retimed_I3833_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3833_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0];
	end
assign N6430 = x_reg_L1_0__retimed_I3833_QOUT;
reg x_reg_L0_23__retimed_I3782_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3782_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650;
	end
assign N6304 = x_reg_L0_23__retimed_I3782_QOUT;
reg x_reg_L0_7__retimed_I3780_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I3780_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912;
	end
assign N6299 = x_reg_L0_7__retimed_I3780_QOUT;
reg x_reg_L1_0__retimed_I3747_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3747_QOUT <= N5654;
	end
assign N6154 = x_reg_L1_0__retimed_I3747_QOUT;
reg x_reg_L1_1__retimed_I3744_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3744_QOUT <= N5647;
	end
assign N6147 = x_reg_L1_1__retimed_I3744_QOUT;
reg x_reg_L1_2__retimed_I3741_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3741_QOUT <= N5640;
	end
assign N6140 = x_reg_L1_2__retimed_I3741_QOUT;
reg x_reg_L1_3__retimed_I3738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3738_QOUT <= N5633;
	end
assign N6133 = x_reg_L1_3__retimed_I3738_QOUT;
reg x_reg_L1_4__retimed_I3735_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3735_QOUT <= N5626;
	end
assign N6126 = x_reg_L1_4__retimed_I3735_QOUT;
reg x_reg_L1_5__retimed_I3732_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3732_QOUT <= N5619;
	end
assign N6119 = x_reg_L1_5__retimed_I3732_QOUT;
reg x_reg_L1_6__retimed_I3729_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3729_QOUT <= N5612;
	end
assign N6112 = x_reg_L1_6__retimed_I3729_QOUT;
reg x_reg_L1_7__retimed_I3726_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3726_QOUT <= N5605;
	end
assign N6105 = x_reg_L1_7__retimed_I3726_QOUT;
reg x_reg_L1_8__retimed_I3723_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3723_QOUT <= N5598;
	end
assign N6098 = x_reg_L1_8__retimed_I3723_QOUT;
reg x_reg_L1_9__retimed_I3720_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I3720_QOUT <= N5591;
	end
assign N6091 = x_reg_L1_9__retimed_I3720_QOUT;
reg x_reg_L1_10__retimed_I3717_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I3717_QOUT <= N5584;
	end
assign N6084 = x_reg_L1_10__retimed_I3717_QOUT;
reg x_reg_L1_11__retimed_I3714_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I3714_QOUT <= N5577;
	end
assign N6077 = x_reg_L1_11__retimed_I3714_QOUT;
reg x_reg_L1_12__retimed_I3711_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3711_QOUT <= N5570;
	end
assign N6070 = x_reg_L1_12__retimed_I3711_QOUT;
reg x_reg_L1_13__retimed_I3708_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3708_QOUT <= N5563;
	end
assign N6063 = x_reg_L1_13__retimed_I3708_QOUT;
reg x_reg_L1_14__retimed_I3705_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I3705_QOUT <= N5556;
	end
assign N6056 = x_reg_L1_14__retimed_I3705_QOUT;
reg x_reg_L1_15__retimed_I3702_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3702_QOUT <= N5549;
	end
assign N6049 = x_reg_L1_15__retimed_I3702_QOUT;
reg x_reg_L1_16__retimed_I3699_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3699_QOUT <= N5542;
	end
assign N6042 = x_reg_L1_16__retimed_I3699_QOUT;
reg x_reg_L1_17__retimed_I3696_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3696_QOUT <= N5535;
	end
assign N6035 = x_reg_L1_17__retimed_I3696_QOUT;
reg x_reg_L1_18__retimed_I3693_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3693_QOUT <= N5528;
	end
assign N6028 = x_reg_L1_18__retimed_I3693_QOUT;
reg x_reg_L1_19__retimed_I3690_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3690_QOUT <= N5521;
	end
assign N6021 = x_reg_L1_19__retimed_I3690_QOUT;
reg x_reg_L1_20__retimed_I3687_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I3687_QOUT <= N5514;
	end
assign N6014 = x_reg_L1_20__retimed_I3687_QOUT;
reg x_reg_L1_21__retimed_I3684_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I3684_QOUT <= N5507;
	end
assign N6007 = x_reg_L1_21__retimed_I3684_QOUT;
reg x_reg_L0_31__retimed_I3681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3681_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6;
	end
assign N6000 = x_reg_L0_31__retimed_I3681_QOUT;
reg x_reg_L0_31__retimed_I3680_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3680_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
	end
assign N5998 = x_reg_L0_31__retimed_I3680_QOUT;
reg x_reg_L0_23__retimed_I3672_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3672_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12;
	end
assign N5974 = x_reg_L0_23__retimed_I3672_QOUT;
reg x_reg_L0_23__retimed_I3671_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3671_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17;
	end
assign N5972 = x_reg_L0_23__retimed_I3671_QOUT;
reg x_reg_L0_22__retimed_I3668_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3668_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
	end
assign N5956 = x_reg_L0_22__retimed_I3668_QOUT;
reg x_reg_L0_31__retimed_I3573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3573_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113;
	end
assign N5720 = x_reg_L0_31__retimed_I3573_QOUT;
reg x_reg_L0_31__retimed_I3572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3572_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122;
	end
assign N5718 = x_reg_L0_31__retimed_I3572_QOUT;
reg x_reg_L0_0__retimed_I3545_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I3545_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0];
	end
assign N5654 = x_reg_L0_0__retimed_I3545_QOUT;
reg x_reg_L0_1__retimed_I3542_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I3542_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1];
	end
assign N5647 = x_reg_L0_1__retimed_I3542_QOUT;
reg x_reg_L0_2__retimed_I3539_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I3539_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2];
	end
assign N5640 = x_reg_L0_2__retimed_I3539_QOUT;
reg x_reg_L0_3__retimed_I3536_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I3536_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3];
	end
assign N5633 = x_reg_L0_3__retimed_I3536_QOUT;
reg x_reg_L0_4__retimed_I3533_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I3533_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4];
	end
assign N5626 = x_reg_L0_4__retimed_I3533_QOUT;
reg x_reg_L0_5__retimed_I3530_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I3530_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5];
	end
assign N5619 = x_reg_L0_5__retimed_I3530_QOUT;
reg x_reg_L0_6__retimed_I3527_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I3527_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6];
	end
assign N5612 = x_reg_L0_6__retimed_I3527_QOUT;
reg x_reg_L0_7__retimed_I3524_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I3524_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7];
	end
assign N5605 = x_reg_L0_7__retimed_I3524_QOUT;
reg x_reg_L0_8__retimed_I3521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I3521_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8];
	end
assign N5598 = x_reg_L0_8__retimed_I3521_QOUT;
reg x_reg_L0_9__retimed_I3518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I3518_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9];
	end
assign N5591 = x_reg_L0_9__retimed_I3518_QOUT;
reg x_reg_L0_10__retimed_I3515_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I3515_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10];
	end
assign N5584 = x_reg_L0_10__retimed_I3515_QOUT;
reg x_reg_L0_11__retimed_I3512_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I3512_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11];
	end
assign N5577 = x_reg_L0_11__retimed_I3512_QOUT;
reg x_reg_L0_12__retimed_I3509_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I3509_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12];
	end
assign N5570 = x_reg_L0_12__retimed_I3509_QOUT;
reg x_reg_L0_13__retimed_I3506_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I3506_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13];
	end
assign N5563 = x_reg_L0_13__retimed_I3506_QOUT;
reg x_reg_L0_14__retimed_I3503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I3503_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14];
	end
assign N5556 = x_reg_L0_14__retimed_I3503_QOUT;
reg x_reg_L0_15__retimed_I3500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I3500_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15];
	end
assign N5549 = x_reg_L0_15__retimed_I3500_QOUT;
reg x_reg_L0_16__retimed_I3497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I3497_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16];
	end
assign N5542 = x_reg_L0_16__retimed_I3497_QOUT;
reg x_reg_L0_17__retimed_I3494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I3494_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17];
	end
assign N5535 = x_reg_L0_17__retimed_I3494_QOUT;
reg x_reg_L0_18__retimed_I3491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I3491_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18];
	end
assign N5528 = x_reg_L0_18__retimed_I3491_QOUT;
reg x_reg_L0_19__retimed_I3488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I3488_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19];
	end
assign N5521 = x_reg_L0_19__retimed_I3488_QOUT;
reg x_reg_L0_20__retimed_I3485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I3485_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20];
	end
assign N5514 = x_reg_L0_20__retimed_I3485_QOUT;
reg x_reg_L0_21__retimed_I3482_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I3482_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21];
	end
assign N5507 = x_reg_L0_21__retimed_I3482_QOUT;
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I0 (.Y(bdw_enable), .A(astall));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083), .A(a_exp[0]), .B(a_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I2 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I3 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194), .A(a_exp[7]), .B(a_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I4 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I5 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I6 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I7 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106), .A(a_man[10]), .B(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I8 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125), .A(a_man[6]), .B(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I9 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114), .A(a_man[8]), .B(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I10 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134), .A(a_man[4]), .B(a_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I11 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I12 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I13 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I14 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I15 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I16 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168), .A(b_exp[0]), .B(b_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I17 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I18 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202), .A(b_exp[7]), .B(b_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I19 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I20 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I21 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I22 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191), .A(b_man[10]), .B(b_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I23 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210), .A(b_man[6]), .B(b_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I24 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199), .A(b_man[8]), .B(b_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I25 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219), .A(b_man[4]), .B(b_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I26 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I27 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I28 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I29 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I30 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I31 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I32 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I33 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I34 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
OR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I35 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I36 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563), .A(b_exp[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I37 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562), .A(b_exp[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I38 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561), .A(b_exp[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I39 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560), .A(b_exp[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I40 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559), .A(b_exp[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I41 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558), .A(b_exp[2]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I42 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557), .A(b_exp[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I43 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556), .A(b_exp[0]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I44 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I45 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I46 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I47 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558), .B(a_exp[2]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I48 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I49 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I50 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561), .B(a_exp[5]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I51 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562), .B(a_exp[6]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I52 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563), .B(a_exp[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I53 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I54 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457), .A(a_man[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I55 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475), .A(b_man[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I56 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544), .A(a_man[21]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I57 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I58 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478), .A(a_man[20]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I59 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I60 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I61 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I62 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410), .A(a_man[19]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I63 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I64 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498), .A(a_man[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I65 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I66 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I67 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431), .A(a_man[17]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I68 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I69 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515), .A(a_man[16]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I70 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I71 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I72 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I73 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489), .A(a_man[11]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I74 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I75 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421), .A(a_man[10]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I76 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I77 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I78 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507), .A(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I79 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I80 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453), .A(a_man[15]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I81 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I82 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535), .A(a_man[14]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I83 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I84 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I85 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468), .A(a_man[13]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I86 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I87 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405), .A(a_man[12]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I88 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I89 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I90 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I91 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444), .A(a_man[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I92 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I93 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I94 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525), .A(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I95 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I96 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461), .A(a_man[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I97 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I98 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I99 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547), .A(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I101 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480), .A(a_man[4]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I104 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I105 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415), .A(a_man[3]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I106 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I107 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501), .A(a_man[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I108 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I109 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I110 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441), .A(b_man[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434), .A(a_man[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434));
OAI31X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I114 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441), .A1(a_man[0]), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I123 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I124 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I125 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I126 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I127 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I128 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I129 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I130 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I131 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I132 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I133 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I134 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I135 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I136 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I137 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I138 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I139 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I140 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I141 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I142 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I143 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I144 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I145 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I146 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I147 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I148 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I149 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I150 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I151 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I152 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I153 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473), .B0(b_man[22]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I154 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I155 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I156 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I157 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I158 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558), .B(a_exp[2]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I159 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I160 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I161 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561), .B(a_exp[5]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I162 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562), .B(a_exp[6]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I163 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572), .A(a_exp[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I164 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I165 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575));
CLKINVX8 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I166 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I167 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I168 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I169 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .A(a_man[7]), .B(b_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I170 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I171 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I172 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I173 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I174 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I175 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I176 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295));
OR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I177 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I178 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I179 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I180 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I181 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I182 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I183 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I184 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I185 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I186 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I187 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I188 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
OAI211X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I189 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I190 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I191 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I192 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I193 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
NOR3BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I194 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]));
NAND2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I195 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I196 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I197 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I198 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556), .B(a_exp[0]));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I199 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I200 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I201 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I202 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I203 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I204 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I205 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I206 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I207 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I208 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I209 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828), .A(b_man[11]), .B(a_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I210 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I211 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I212 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I213 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I214 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I215 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I216 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I217 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835), .A(b_man[14]), .B(a_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I218 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I219 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842), .A(b_man[13]), .B(a_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I220 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I221 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I222 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I223 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I224 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I225 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I226 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I227 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I228 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .A(b_man[20]), .B(a_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I229 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .A(b_man[19]), .B(a_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I230 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I231 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I232 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I233 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I234 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I235 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I236 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I237 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I238 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I239 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I240 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I241 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I242 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I243 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I244 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I245 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I246 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I247 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I248 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I249 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .A(a_man[6]), .B(b_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I250 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I251 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I252 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I253 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I254 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I255 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I256 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I257 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I258 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I259 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I260 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I261 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I262 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I263 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I264 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I265 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I266 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I267 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I269 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I270 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I271 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I272 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I273 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I274 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I275 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I276 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I277 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I278 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I279 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I280 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I281 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I282 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I283 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I284 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I285 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I286 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I287 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I288 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I289 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629), .A(a_man[5]), .B(b_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I290 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I291 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I292 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I293 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613), .A(a_man[4]), .B(b_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I294 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I295 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I296 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058), .A(b_man[4]), .B(a_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I297 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I298 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I299 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I300 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I301 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I302 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I303 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I304 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I305 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I306 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I307 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I308 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I309 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I310 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I311 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I312 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849), .A(b_man[3]), .B(a_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I313 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I314 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I315 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I316 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I317 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I318 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I319 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I320 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I321 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I322 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I323 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I324 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .A(a_man[3]), .B(b_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I325 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I326 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I327 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I328 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I329 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I330 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I331 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I332 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I333 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I334 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I335 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I336 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I337 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I338 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I339 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I340 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I341 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385));
OR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I342 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I343 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366), .A(a_man[1]), .B(b_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I344 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I345 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I346 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I347 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I348 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I349 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I350 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I351 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I352 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I353 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I354 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I355 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I356 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I357 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I358 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I359 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .A(a_man[0]), .B(b_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I360 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I361 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I362 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .A(b_man[0]), .B(a_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I363 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I364 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I365 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I366 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I367 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I368 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I369 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I370 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I371 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I372 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]));
XOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I373 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I374 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I375 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I376 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I377 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I378 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I379 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I380 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I381 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I382 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I383 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I384 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I385 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I386 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I387 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I388 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I390 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I391 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I392 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I393 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I394 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I396 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I397 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I398 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I399 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I400 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I401 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I402 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I403 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I404 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I407 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I409 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I412 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I413 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I415 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I416 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I417 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I418 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I419 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I420 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I421 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I422 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I423 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I424 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I425 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I427 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I428 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I429 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I430 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I431 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I432 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I433 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I434 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I435 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I436 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I437 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I438 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I439 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I440 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I441 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I442 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I443 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I444 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I445 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I446 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I447 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I448 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I449 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I450 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I451 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I452 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I453 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I454 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I455 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I456 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332));
AOI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I457 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I458 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I459 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I460 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I461 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I462 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I463 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I464 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I465 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I466 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I467 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I468 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I469 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I470 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I471 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635), .A(N10166), .B(N10168));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I472 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601), .AN(N9398), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I473 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606), .A(N9576), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I474 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I475 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I476 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718), .A0N(N9382), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643), .B0(N9565));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I477 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I478 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709), .A0N(N9374), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718), .B0(N9557));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I479 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I480 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .A(a_man[8]), .B(b_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I481 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I482 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I483 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I484 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I485 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I486 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709), .B(N9366));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I487 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718), .B(N9374));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I488 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I489 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643), .B(N9382));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I490 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611), .A(N10168));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I491 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635), .A0N(N9431), .A1N(N9433), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I492 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635), .B(N9398));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I493 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I494 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864));
INVXL buf1_A_I5405 (.Y(N10666), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599));
INVXL buf1_A_I5406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667), .A(N10666));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I496 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691), .A0N(N9406), .A1N(N9404), .B0(N9422));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I497 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691), .B(N9390));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I498 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .A(N9404), .B(N9406));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I499 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I500 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I501 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I502 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I503 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .A(N10157), .B(N10159));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I504 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I505 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I506 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I507 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I508 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I509 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I510 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I511 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .B(N8521));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I512 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I513 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I514 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I515 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .A(a_man[15]), .B(b_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I516 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I517 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I518 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I519 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I520 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I521 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .A(a_man[14]), .B(b_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I522 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I523 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I524 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I525 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I526 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I527 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .A(a_man[13]), .B(b_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I528 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I529 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I530 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I531 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I532 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I533 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .A(a_man[12]), .B(b_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I534 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I535 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I536 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I537 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I538 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I539 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .A(a_man[11]), .B(b_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I540 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I541 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I542 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I543 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I544 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I545 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .A(a_man[10]), .B(b_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I546 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I547 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I548 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I549 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I550 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I551 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .A(a_man[9]), .B(b_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I552 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I553 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I554 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I555 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I556 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I557 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I558 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612), .A0N(N9366), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709), .B0(N9549));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I559 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I560 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583), .A0N(N9358), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612), .B0(N9541));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I561 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I562 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616), .A0N(N9350), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583), .B0(N9533));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I563 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I564 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717), .A0N(N9342), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616), .B0(N9525));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I565 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I566 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .A0N(N9334), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717), .B0(N9517));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I567 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I568 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664), .A0N(N9326), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .B0(N9509));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I569 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I570 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659), .A0N(N9318), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664), .B0(N9501));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I571 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I572 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723), .A0N(N9310), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659), .B0(N9493));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I573 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .A(a_man[16]), .B(b_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I574 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I575 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I576 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I577 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723), .B(N9302));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I578 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659), .B(N9310));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I579 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I580 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664), .B(N9318));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I581 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .B(N9326));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I582 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I583 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I584 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717), .B(N9334));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I585 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616), .B(N9342));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I586 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I587 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583), .B(N9350));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I588 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612), .B(N9358));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I589 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I590 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I591 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I592 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I593 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .A(a_man[19]), .B(b_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I594 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I595 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I596 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I597 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .A(a_man[18]), .B(b_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I598 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I599 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I600 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I601 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I602 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .A(a_man[17]), .B(b_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I603 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I604 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I605 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I606 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I607 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I608 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699), .A0N(N9302), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723), .B0(N9485));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I609 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I610 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .A0N(N9295), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699), .B0(N9477));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I611 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I612 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701), .A0N(N9288), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .B0(N9469));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I613 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I614 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578), .A0N(N9281), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701), .B0(N9461));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I615 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .A(a_man[20]), .B(b_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I616 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I617 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I618 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I619 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578), .B(N9274));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I620 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701), .B(N9281));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I621 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I622 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .B(N9288));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I623 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699), .B(N9295));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I624 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I625 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I626 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .A(a_man[21]), .B(b_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I627 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I628 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I629 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I630 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I631 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666), .A0N(N9274), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578), .B0(N9453));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I632 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I633 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672), .A0N(N9267), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666), .B0(N9445));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I634 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .A(a_man[22]), .B(b_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I635 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I636 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I637 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I638 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672), .B(N9260));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I639 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666), .B(N9267));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I640 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I641 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I642 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I643 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I644 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594), .A0N(N9260), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672), .B0(N9437));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I645 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624), .A(N9246), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I646 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]), .A(N9251), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I647 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594), .B(N9246));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I648 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I649 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I650 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I651 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I652 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I653 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I654 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893));
OA21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I655 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I656 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I657 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I658 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I659 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I660 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I661 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729), .A(N7068), .B(N7070));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I662 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I663 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I664 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I665 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I666 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I667 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I668 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I669 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I670 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I671 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I672 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
BUFX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I673 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I674 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I675 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I676 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I677 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I678 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I679 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869), .AN(N8521), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I680 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I681 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I682 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I683 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I684 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I685 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I686 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831), .A1(N8990), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I687 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I688 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I689 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I690 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4860), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I691 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4881), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I692 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4902), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4860), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4881));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I693 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4877), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4902));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I694 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4889), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I695 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I696 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4838), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4889), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I697 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4824), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I698 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4847), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I699 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4866), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4847));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I700 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4917), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4838), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4866));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I701 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4877), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4917));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I702 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I703 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I704 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I705 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
BUFX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I706 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I707 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I708 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I709 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I710 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870), .A(N8941), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831));
NAND2BX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I711 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I712 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I713 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4901), .AN(N8941), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I714 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4828), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892));
AO21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I715 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4828));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I716 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I717 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I718 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I719 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I720 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I721 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I722 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285), .A(N8521), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I723 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I724 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I725 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I726 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I727 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I728 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I729 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I730 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I731 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I732 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I733 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I734 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I735 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5284), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I736 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214), .A(N8528), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I737 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I738 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I739 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143), .A(N8536), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I740 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I741 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I742 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I743 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I744 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I745 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I746 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I747 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I748 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I749 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I750 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I751 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I752 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5284), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I753 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I754 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223), .A(N8536), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I755 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I756 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I757 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I758 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5157), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I759 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I760 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I761 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I762 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5157), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I763 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I764 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I765 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I766 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I767 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I768 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I769 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I770 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I771 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I772 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I773 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I774 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I775 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I776 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I777 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I778 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I779 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I780 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I781 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I782 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I783 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I784 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I785 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I786 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I787 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I788 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I789 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I790 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128), .A(N8521), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I791 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I792 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I793 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I794 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I795 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I796 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258), .A(N8528), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I797 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I798 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I799 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I800 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I801 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I802 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I803 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I804 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I805 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I806 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I807 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I808 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I809 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I810 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I811 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I812 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I813 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I814 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I815 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I816 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I817 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I818 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I819 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I820 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I821 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I822 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I823 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I824 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I825 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I826 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I827 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I828 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I829 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I830 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I831 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I832 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I833 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I834 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I835 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I836 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I837 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I838 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I839 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I840 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5576), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I841 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I842 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I843 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I844 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I845 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I846 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I847 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I848 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I849 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I850 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I851 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I852 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I853 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I854 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I855 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I856 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I857 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I858 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I859 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I860 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I861 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I862 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48), .A(b_sign), .B(a_sign), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I863 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I864 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I865 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I866 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I867 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I868 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I869 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30));
AO21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I870 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I871 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I872 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I873 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I874 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I875 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631), .A(N8578), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I876 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631), .B(N8480), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I877 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280), .A(N8017), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I878 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I879 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I880 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]), .B(N8110), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I881 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I882 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I883 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I884 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I885 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633), .A(N8203), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632));
NOR4X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I886 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269), .A(N8100), .B(N8102), .C(N8104), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I887 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I888 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I889 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I890 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314));
NAND4X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I891 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I892 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072));
CLKAND2X3 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I893 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5576), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
NAND4X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I894 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8080), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I895 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8080));
NAND3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I896 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8086), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I897 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8086));
NAND3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I898 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8139), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I899 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8139));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I900 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13744), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]), .A(N7272), .B(N7270), .CI(N10193));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I901 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13695), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .A(N7259), .B(N7257), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13744));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I902 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13732), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .A(N7241), .B(N7239), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I903 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I904 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I905 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754), .A(N10123), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I906 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724), .A(N10111), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I907 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13685), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]), .A(N7223), .B(N7221), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13732));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I908 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13722), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .A(N7205), .B(N7203), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13685));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I909 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I910 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I911 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13746), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .A(N7187), .B(N7185), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13722));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I912 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]), .A(b_exp[6]), .B(a_exp[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I913 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I914 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]), .A(N7169), .B(N7167), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13746));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I915 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13719), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]));
OR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I916 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13692), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I917 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]), .A(b_exp[7]), .B(a_exp[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I918 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742), .A(N10116));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I919 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446), .A(N10116));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I920 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686), .A(N7151), .B(N7149), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I921 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I5377 (.Y(N10610), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I5378 (.Y(N10611), .A(N10610));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I922 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683), .A(N7091), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I923 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I924 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13730), .A(N7091), .B(N10611));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I925 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13699), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686));
NAND3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I926 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13699), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13738), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13730));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I927 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I928 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I929 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I930 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I931 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I932 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707));
AO21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I933 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642), .A0(N7501), .A1(N10193), .B0(N7505));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I934 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754), .A(N7427), .B(N7429), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I935 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .A(N7099), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I936 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13740), .A(N7083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I937 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13701), .A(N7038), .B(N7040), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13740));
OAI31X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I938 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__71), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13719), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13692), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13706), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13701));
INVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I939 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__71));
INVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I940 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875));
INVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I941 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
NOR2BX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I942 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .AN(N6655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I943 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893), .A(rm[0]), .B(rm[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I944 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7), .A(rm[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I945 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I946 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I947 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I948 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .B(N6837));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I949 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .A(N6655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I950 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I951 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I952 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]), .A(N7661), .B(N7663));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I953 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I954 (.Y(x[22]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I955 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I956 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[21]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[21]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I957 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]), .A(N7931), .B(N7933));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I958 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I959 (.Y(x[21]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6007), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I960 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[20]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[20]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I961 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I962 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I963 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(N10173));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I964 (.Y(x[20]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6014), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I965 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[19]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[19]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I966 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I967 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(N6601));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I968 (.Y(x[19]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6021), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I969 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[18]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[18]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I970 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I971 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I972 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I973 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(N6592));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I974 (.Y(x[18]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6028), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I975 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[17]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[17]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I976 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I977 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I978 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(N6583));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I979 (.Y(x[17]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6035), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I980 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[16]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[16]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I981 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I982 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I983 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(N6574));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I984 (.Y(x[16]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I985 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[15]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[15]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I986 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I987 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(N6565));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I988 (.Y(x[15]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6049), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I989 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[14]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[14]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I990 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I991 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I992 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I993 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I994 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I995 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I996 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I997 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I998 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I999 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1000 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1001 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1002 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(N10175));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1003 (.Y(x[14]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6056), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1004 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[13]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[13]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1005 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1006 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(N6547));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1007 (.Y(x[13]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6063), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1008 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[12]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1009 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1010 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1011 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1012 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(N6538));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1013 (.Y(x[12]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6070), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1014 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[11]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[11]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1015 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1016 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(N6529));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1017 (.Y(x[11]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6077), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1018 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[10]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[10]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1019 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1020 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1021 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1022 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(N6520));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1023 (.Y(x[10]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6084), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1024 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[9]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[9]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1025 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1026 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(N6511));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1027 (.Y(x[9]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6091), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1028 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[8]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1029 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1030 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1031 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(N6502));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1032 (.Y(x[8]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6098), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1033 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[7]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[7]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1034 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1035 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6493));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1036 (.Y(x[7]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6105), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1037 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[6]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[6]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1038 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1039 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1040 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1041 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6484));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1042 (.Y(x[6]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6112), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1043 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[5]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[5]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1044 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1045 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6475));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1046 (.Y(x[5]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6119), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1047 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[4]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1048 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1049 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1050 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6466));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1051 (.Y(x[4]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6126), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1052 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[3]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[3]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1053 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1054 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6457));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1055 (.Y(x[3]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6133), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1056 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[2]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1057 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1058 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1059 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1060 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1061 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1062 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1063 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6448));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1064 (.Y(x[2]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6140), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1065 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[1]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1066 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1067 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6439));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1068 (.Y(x[1]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6147), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1069 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[0]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[0]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1070 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1071 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(N6430));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1072 (.Y(x[0]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N6154), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926));
INVXL buf1_A_I5407 (.Y(N10671), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686));
INVXL buf1_A_I5408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]), .A(N10671));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1074 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .A(N6673), .B(N6671), .C(N6655), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1075 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1076 (.Y(x[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1077 (.Y(x[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1078 (.Y(x[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1079 (.Y(x[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1080 (.Y(x[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1081 (.Y(x[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1082 (.Y(x[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1083 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1084 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651), .A(N6842), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1085 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]), .A(N6671), .B(N6673), .C(N6655), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1086 (.Y(x[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1087 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881), .A(a_sign), .B(b_sign));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1088 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1089 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1090 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064), .A0(a_sign), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_sign));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1091 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1092 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1093 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116), .A(N5998), .B(N6000), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1094 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_5_I1095 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[31]), .A(N5720), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116), .S0(N5718));
reg x_reg_L1_31__I1159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I1159_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[31];
	end
assign x[31] = x_reg_L1_31__I1159_QOUT;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[0] = x[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[1] = x[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[2] = x[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[3] = x[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[4] = x[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[5] = x[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[6] = x[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[7] = x[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[8] = x[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[9] = x[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[10] = x[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[11] = x[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[12] = x[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[13] = x[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[14] = x[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[15] = x[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[16] = x[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[17] = x[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[18] = x[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[19] = x[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[20] = x[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[21] = x[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[22] = x[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[23] = x[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[24] = x[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[25] = x[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[26] = x[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[27] = x[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[28] = x[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[29] = x[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[30] = x[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[28] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  v7XzSw3cohw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



