/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:25:11 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__53,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4799,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4818,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4865,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4898,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5201,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5237,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5244,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5249,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5259,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5345,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6158,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6187,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6200,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6207,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6226,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6239,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6244,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6249,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6256,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6262,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6288,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6292,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6303,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6311,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6315,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6334,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6393,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6395,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6440,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6476,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6764,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6818,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6987,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7209,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7216,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7255,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7292,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7304,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7345,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7625,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7640,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7737,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7755,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7791,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7941,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7976,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8067,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8100,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8112,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8118,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8276,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8435,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8440,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17458,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17463,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17590,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17637,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17818,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17979;
wire N6622,N6624,N6662,N6666,N6673,N6680,N6687 
	,N6694,N6701,N6708,N6715,N6722,N6729,N6732,N6739 
	,N6746,N6753,N6760,N6767,N6774,N6781,N6788,N6795 
	,N6802,N6809,N6821,N6955,N6957,N6959,N6992,N6997 
	,N6999,N7090,N7208,N7210,N7317,N7325,N7327,N7354 
	,N7356,N7358,N7364,N7472,N7476,N7682,N7705,N7713 
	,N7719,N7727,N7735,N8267,N8274,N8454,N8457,N8467 
	,N8469,N8472,N8621,N8625,N8641,N8643,N8650,N8652 
	,N8657,N8662,N8664,N8667,N8669,N8671,N8678,N8683 
	,N8685,N8690,N8692,N8696,N8698,N8700,N8703,N8707 
	,N8714,N8721,N8726,N8728,N8733,N8735,N8738,N8742 
	,N8749,N8756,N8761,N8770,N8773,N8775,N8785,N8803 
	,N8812,N8835,N8981,N9037,N9662,N9663,N9664,N9665 
	,N9666,N9667,N9668,N9669,N9670,N9671,N9672,N9673 
	,N9718,N9719,N9720,N9721;
reg x_reg_24__retimed_I5353_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5353_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[0];
	end
assign N9037 = x_reg_24__retimed_I5353_QOUT;
reg x_reg_24__retimed_I5326_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5326_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653;
	end
assign N8981 = x_reg_24__retimed_I5326_QOUT;
reg x_reg_24__retimed_I5301_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5301_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17637;
	end
assign N8835 = x_reg_24__retimed_I5301_QOUT;
reg x_reg_24__retimed_I5292_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5292_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7603;
	end
assign N8812 = x_reg_24__retimed_I5292_QOUT;
reg x_reg_24__retimed_I5289_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5289_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734;
	end
assign N8803 = x_reg_24__retimed_I5289_QOUT;
reg x_reg_24__retimed_I5283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5283_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5];
	end
assign N8785 = x_reg_24__retimed_I5283_QOUT;
reg x_reg_24__retimed_I5280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5280_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10721;
	end
assign N8775 = x_reg_24__retimed_I5280_QOUT;
reg x_reg_24__retimed_I5279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5279_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10715;
	end
assign N8773 = x_reg_24__retimed_I5279_QOUT;
reg x_reg_24__retimed_I5278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5278_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17];
	end
assign N8770 = x_reg_24__retimed_I5278_QOUT;
reg x_reg_24__retimed_I5274_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5274_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16];
	end
assign N8761 = x_reg_24__retimed_I5274_QOUT;
reg x_reg_24__retimed_I5272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5272_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22];
	end
assign N8756 = x_reg_24__retimed_I5272_QOUT;
reg x_reg_24__retimed_I5269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5269_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21];
	end
assign N8749 = x_reg_24__retimed_I5269_QOUT;
reg x_reg_24__retimed_I5266_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5266_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23];
	end
assign N8742 = x_reg_24__retimed_I5266_QOUT;
reg x_reg_24__retimed_I5264_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5264_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738;
	end
assign N8738 = x_reg_24__retimed_I5264_QOUT;
reg x_reg_24__retimed_I5263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5263_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9];
	end
assign N8735 = x_reg_24__retimed_I5263_QOUT;
reg x_reg_24__retimed_I5262_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5262_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1];
	end
assign N8733 = x_reg_24__retimed_I5262_QOUT;
reg x_reg_24__retimed_I5260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5260_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15];
	end
assign N8728 = x_reg_24__retimed_I5260_QOUT;
reg x_reg_24__retimed_I5259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5259_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7];
	end
assign N8726 = x_reg_24__retimed_I5259_QOUT;
reg x_reg_24__retimed_I5257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5257_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20];
	end
assign N8721 = x_reg_24__retimed_I5257_QOUT;
reg x_reg_24__retimed_I5254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5254_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19];
	end
assign N8714 = x_reg_24__retimed_I5254_QOUT;
reg x_reg_24__retimed_I5251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5251_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18];
	end
assign N8707 = x_reg_24__retimed_I5251_QOUT;
reg x_reg_24__retimed_I5249_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5249_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737;
	end
assign N8703 = x_reg_24__retimed_I5249_QOUT;
reg x_reg_24__retimed_I5248_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5248_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8];
	end
assign N8700 = x_reg_24__retimed_I5248_QOUT;
reg x_reg_24__retimed_I5247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5247_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0];
	end
assign N8698 = x_reg_24__retimed_I5247_QOUT;
reg x_reg_24__retimed_I5246_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5246_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735;
	end
assign N8696 = x_reg_24__retimed_I5246_QOUT;
reg x_reg_24__retimed_I5245_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5245_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10];
	end
assign N8692 = x_reg_24__retimed_I5245_QOUT;
reg x_reg_24__retimed_I5244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5244_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2];
	end
assign N8690 = x_reg_24__retimed_I5244_QOUT;
reg x_reg_24__retimed_I5242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5242_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11];
	end
assign N8685 = x_reg_24__retimed_I5242_QOUT;
reg x_reg_24__retimed_I5241_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5241_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3];
	end
assign N8683 = x_reg_24__retimed_I5241_QOUT;
reg x_reg_24__retimed_I5239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5239_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13];
	end
assign N8678 = x_reg_24__retimed_I5239_QOUT;
reg x_reg_24__retimed_I5236_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5236_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12];
	end
assign N8671 = x_reg_24__retimed_I5236_QOUT;
reg x_reg_24__retimed_I5235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5235_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4];
	end
assign N8669 = x_reg_24__retimed_I5235_QOUT;
reg x_reg_24__retimed_I5234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5234_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736;
	end
assign N8667 = x_reg_24__retimed_I5234_QOUT;
reg x_reg_24__retimed_I5233_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5233_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14];
	end
assign N8664 = x_reg_24__retimed_I5233_QOUT;
reg x_reg_24__retimed_I5232_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5232_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6];
	end
assign N8662 = x_reg_24__retimed_I5232_QOUT;
reg x_reg_24__retimed_I5230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5230_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17626;
	end
assign N8657 = x_reg_24__retimed_I5230_QOUT;
reg x_reg_24__retimed_I5228_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5228_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17638;
	end
assign N8652 = x_reg_24__retimed_I5228_QOUT;
reg x_reg_24__retimed_I5227_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5227_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17628;
	end
assign N8650 = x_reg_24__retimed_I5227_QOUT;
reg x_reg_24__retimed_I5224_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5224_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17664;
	end
assign N8643 = x_reg_24__retimed_I5224_QOUT;
reg x_reg_24__retimed_I5223_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5223_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663;
	end
assign N8641 = x_reg_24__retimed_I5223_QOUT;
reg x_reg_24__retimed_I5217_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5217_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693;
	end
assign N8625 = x_reg_24__retimed_I5217_QOUT;
reg x_reg_24__retimed_I5215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5215_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[1];
	end
assign N8621 = x_reg_24__retimed_I5215_QOUT;
reg x_reg_24__retimed_I5160_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5160_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620;
	end
assign N8472 = x_reg_24__retimed_I5160_QOUT;
reg x_reg_24__retimed_I5159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5159_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234;
	end
assign N8469 = x_reg_24__retimed_I5159_QOUT;
assign N9662 = !N8469;
assign N9663 = !N9662;
assign N9664 = !N8469;
assign N9718 = !N9664;
assign N9719 = !N9718;
assign N9720 = !N9664;
assign N9721 = !N9720;
assign N9669 = !N9721;
assign N9668 = !N9719;
assign N9667 = !N9721;
assign N9666 = !N9721;
assign N9665 = !N9721;
reg x_reg_24__retimed_I5158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5158_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7211;
	end
assign N8467 = x_reg_24__retimed_I5158_QOUT;
reg x_reg_24__retimed_I5154_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5154_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4;
	end
assign N8457 = x_reg_24__retimed_I5154_QOUT;
reg x_reg_24__retimed_I5153_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5153_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43;
	end
assign N8454 = x_reg_24__retimed_I5153_QOUT;
reg x_reg_24__retimed_I5085_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5085_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635;
	end
assign N8274 = x_reg_24__retimed_I5085_QOUT;
reg x_reg_24__retimed_I5082_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I5082_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7640;
	end
assign N8267 = x_reg_24__retimed_I5082_QOUT;
reg x_reg_24__retimed_I4896_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4896_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[3];
	end
assign N7735 = x_reg_24__retimed_I4896_QOUT;
reg x_reg_24__retimed_I4894_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4894_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[4];
	end
assign N7727 = x_reg_24__retimed_I4894_QOUT;
reg x_reg_24__retimed_I4892_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4892_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[1];
	end
assign N7719 = x_reg_24__retimed_I4892_QOUT;
reg x_reg_24__retimed_I4890_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4890_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[2];
	end
assign N7713 = x_reg_24__retimed_I4890_QOUT;
reg x_reg_24__retimed_I4888_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4888_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[0];
	end
assign N7705 = x_reg_24__retimed_I4888_QOUT;
reg x_reg_24__retimed_I4881_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4881_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045;
	end
assign N7682 = x_reg_24__retimed_I4881_QOUT;
reg x_reg_24__retimed_I4811_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4811_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24];
	end
assign N7476 = x_reg_24__retimed_I4811_QOUT;
reg x_reg_24__retimed_I4809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4809_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25];
	end
assign N7472 = x_reg_24__retimed_I4809_QOUT;
reg x_reg_24__retimed_I4773_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4773_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8015;
	end
assign N7364 = x_reg_24__retimed_I4773_QOUT;
reg x_reg_24__retimed_I4772_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4772_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8058;
	end
assign N7358 = x_reg_24__retimed_I4772_QOUT;
reg x_reg_24__retimed_I4771_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4771_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056;
	end
assign N7356 = x_reg_24__retimed_I4771_QOUT;
reg x_reg_24__retimed_I4770_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4770_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042;
	end
assign N7354 = x_reg_24__retimed_I4770_QOUT;
reg x_reg_24__retimed_I4760_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4760_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8037;
	end
assign N7327 = x_reg_24__retimed_I4760_QOUT;
reg x_reg_24__retimed_I4759_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4759_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8057;
	end
assign N7325 = x_reg_24__retimed_I4759_QOUT;
reg x_reg_24__retimed_I4756_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4756_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8111;
	end
assign N7317 = x_reg_24__retimed_I4756_QOUT;
reg x_reg_24__retimed_I4720_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4720_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8112;
	end
assign N7210 = x_reg_24__retimed_I4720_QOUT;
reg x_reg_24__retimed_I4719_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4719_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8094;
	end
assign N7208 = x_reg_24__retimed_I4719_QOUT;
reg x_reg_24__retimed_I4676_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__retimed_I4676_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17483;
	end
assign N7090 = x_reg_24__retimed_I4676_QOUT;
reg x_reg_23__retimed_I4639_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I4639_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8243;
	end
assign N6999 = x_reg_23__retimed_I4639_QOUT;
reg x_reg_23__retimed_I4638_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I4638_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634;
	end
assign N6997 = x_reg_23__retimed_I4638_QOUT;
reg x_reg_22__retimed_I4636_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4636_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8339;
	end
assign N6992 = x_reg_22__retimed_I4636_QOUT;
reg x_reg_31__retimed_I4632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I4632_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[5];
	end
assign N6959 = x_reg_31__retimed_I4632_QOUT;
reg x_reg_31__retimed_I4631_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I4631_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48;
	end
assign N6957 = x_reg_31__retimed_I4631_QOUT;
reg x_reg_31__retimed_I4630_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I4630_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6;
	end
assign N6955 = x_reg_31__retimed_I4630_QOUT;
reg x_reg_23__retimed_I4579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I4579_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8253;
	end
assign N6821 = x_reg_23__retimed_I4579_QOUT;
reg x_reg_21__retimed_I4574_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I4574_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[21];
	end
assign N6809 = x_reg_21__retimed_I4574_QOUT;
reg x_reg_20__retimed_I4571_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I4571_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[20];
	end
assign N6802 = x_reg_20__retimed_I4571_QOUT;
reg x_reg_17__retimed_I4568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I4568_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[17];
	end
assign N6795 = x_reg_17__retimed_I4568_QOUT;
reg x_reg_13__retimed_I4565_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I4565_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[13];
	end
assign N6788 = x_reg_13__retimed_I4565_QOUT;
reg x_reg_12__retimed_I4562_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I4562_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[12];
	end
assign N6781 = x_reg_12__retimed_I4562_QOUT;
reg x_reg_11__retimed_I4559_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I4559_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[11];
	end
assign N6774 = x_reg_11__retimed_I4559_QOUT;
reg x_reg_10__retimed_I4556_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I4556_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[10];
	end
assign N6767 = x_reg_10__retimed_I4556_QOUT;
reg x_reg_8__retimed_I4553_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I4553_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[8];
	end
assign N6760 = x_reg_8__retimed_I4553_QOUT;
reg x_reg_6__retimed_I4550_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I4550_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[6];
	end
assign N6753 = x_reg_6__retimed_I4550_QOUT;
reg x_reg_3__retimed_I4547_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I4547_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[3];
	end
assign N6746 = x_reg_3__retimed_I4547_QOUT;
reg x_reg_2__retimed_I4544_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I4544_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[2];
	end
assign N6739 = x_reg_2__retimed_I4544_QOUT;
reg x_reg_0__retimed_I4541_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I4541_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[0];
	end
assign N6732 = x_reg_0__retimed_I4541_QOUT;
reg x_reg_19__retimed_I4540_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I4540_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[19];
	end
assign N6729 = x_reg_19__retimed_I4540_QOUT;
reg x_reg_18__retimed_I4537_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I4537_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[18];
	end
assign N6722 = x_reg_18__retimed_I4537_QOUT;
reg x_reg_16__retimed_I4534_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I4534_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[16];
	end
assign N6715 = x_reg_16__retimed_I4534_QOUT;
reg x_reg_15__retimed_I4531_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4531_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[15];
	end
assign N6708 = x_reg_15__retimed_I4531_QOUT;
reg x_reg_14__retimed_I4528_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I4528_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[14];
	end
assign N6701 = x_reg_14__retimed_I4528_QOUT;
reg x_reg_9__retimed_I4525_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I4525_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[9];
	end
assign N6694 = x_reg_9__retimed_I4525_QOUT;
reg x_reg_7__retimed_I4522_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I4522_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[7];
	end
assign N6687 = x_reg_7__retimed_I4522_QOUT;
reg x_reg_5__retimed_I4519_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I4519_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[5];
	end
assign N6680 = x_reg_5__retimed_I4519_QOUT;
reg x_reg_4__retimed_I4516_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I4516_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[4];
	end
assign N6673 = x_reg_4__retimed_I4516_QOUT;
reg x_reg_1__retimed_I4513_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I4513_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[1];
	end
assign N6666 = x_reg_1__retimed_I4513_QOUT;
reg x_reg_1__retimed_I4511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I4511_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63;
	end
assign N6662 = x_reg_1__retimed_I4511_QOUT;
assign N9670 = !N6662;
assign N9671 = !N9670;
assign N9672 = !N6662;
assign N9673 = !N9672;
reg x_reg_31__retimed_I4508_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I4508_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7191;
	end
assign N6624 = x_reg_31__retimed_I4508_QOUT;
reg x_reg_31__retimed_I4507_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I4507_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7182;
	end
assign N6622 = x_reg_31__retimed_I4507_QOUT;
assign bdw_enable = !astall;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643 = !a_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563 = !b_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682 = !(a_exp[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562 = !b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635 = !(a_exp[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561 = !b_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697 = !(a_exp[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560 = !b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650 = !(a_exp[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559 = !b_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602 = !(a_exp[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558 = !b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666 = !(a_exp[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557 = !b_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614 = !(a_exp[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556 = !b_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17569 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594 = !(a_exp[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640 = !(a_exp[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687 = !(a_exp[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625 = !(a_exp[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674 = !(a_exp[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609 = !(a_exp[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659 = !(a_exp[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4603 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4603);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17576 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17590 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17569 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17576);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677 = !(a_exp[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843 = !a_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861 = b_man[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864 = !a_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4865 = !(b_man[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931 = !a_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812 = !(b_man[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4891 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4865 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4891);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796 = !a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917 = !(b_man[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884 = !a_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4819 = !(b_man[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4819);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817 = !a_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871 = !(b_man[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901 = !a_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4924 = !(b_man[16] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4873 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4924);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17571 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4873 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922 = !a_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4878 = !(b_man[14] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839 = !a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825 = !(b_man[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4878 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791 = !a_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4832 = !(b_man[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854 = !a_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929 = !(b_man[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4853 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4832 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4853);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829 = !a_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4889 = !(b_man[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893 = !a_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837 = !(b_man[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4836 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4889 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807 = !a_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875 = !a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882 = !(b_man[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807) & (!b_man[10])) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4824 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4836 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4938 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4824);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847 = !a_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4841 = !(b_man[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912 = !a_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790 = !(b_man[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4841 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934 = !a_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892 = !(b_man[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866 = !a_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4794 = !(b_man[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4814 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4794);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4890 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4814);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338 = !a_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4898 = !(b_man[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801 = !a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846 = !(b_man[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4881 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4898 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911 = !b_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820 = !a_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4800 = !(b_man[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4835 = !(b_man[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4914 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911 | a_man[0]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4800) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4835);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4933 = !(b_man[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4880 = !(b_man[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4848 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4933)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4880);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4923 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4881) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4848);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4828 = !(b_man[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4927 = !(b_man[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4935 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4828)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4927);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4874 = !(b_man[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4823 = !(b_man[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4868 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4874) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4823);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4856 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4935 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4868);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4818 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4923) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4890)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4856);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4921 = !(b_man[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4869 = !(b_man[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4802 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4921)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4869);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4816 = !(b_man[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4915 = !(b_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4888 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4816) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4915);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4792 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4802) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4888);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4863 = !(b_man[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4810 = !(b_man[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4822 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4863) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4810);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4910 = !(b_man[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4857 = !(b_man[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4906 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4910)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4857);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4876 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4822 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4906);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4903 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4792) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4876);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17578 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4818 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4938) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4903);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4805 = !(b_man[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4904 = !(b_man[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4840 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4805) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4904);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4851 = !(b_man[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4799 = !(b_man[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4926 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4851) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4799);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4809 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4926);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4897 = !(b_man[20] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4845 = !(b_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4859 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4897)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4845);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4830 = b_man[22] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4894 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4859 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4830);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17586 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4809) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4894));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17595 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17578) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17571)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17586);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17580 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17595);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17590 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17580);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6017 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6017;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25] = a_sign ^ b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[2] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N567 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N567) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N566 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N566) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5114 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17869 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17859 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17859) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17869));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4611 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4611) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N569 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N569) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5119 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4668 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4668);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4649 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5094 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4649) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4665 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N572 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4665 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N572) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5094);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4601 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4601) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4613 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N571 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4613 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N571) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4664 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4664) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4676 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N570 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4676 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N570) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5123 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5119) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5114)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5123);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17818 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17825 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17818 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17825);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17830 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17805 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17830 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17805);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17391 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17391);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5233 = !b_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[40] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5233));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5206 = !b_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[39] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5206));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N565 = (!a_exp[0]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N565) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[39]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5249 = !b_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[36] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5249));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5222 = !b_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[35] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5222));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[35]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5164 = !b_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[42] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5164));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5259 = !b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[41] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5259));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[41]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[42]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5180 = !b_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[38] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5180));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5153 = !b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[37] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5153));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[37]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5141 = !b_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5141));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5237 = !b_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5237));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[31]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433 = !b_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5253 = !b_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5253));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[27]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5195 = !b_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[34] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5195));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5168 = !b_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5168));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[33]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5210 = !b_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5210));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5184 = !b_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5184));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[29]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5201 = !b_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[48] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5201));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5175 = !b_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[47] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5175));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[47]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[48]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5217 = !b_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[44] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5217));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5191 = !b_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[43] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[43]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5148 = !b_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[46] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5148));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5244 = !b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[45] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5244));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[45]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[46]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[27] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6374 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[38]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[34]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[40]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[36]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[30]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224 = !a_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[26]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[32]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[28]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[46]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[47]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[42]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[48]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[44]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[45]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10782 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[26]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10782;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[26]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17372 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17371 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17372);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17371 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[2] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[5] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5922 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[8] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5901 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5899 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5922 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5901);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17814 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5899);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[10] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5931 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[10] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5518 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5518));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5919 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17808 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5931 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5919;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17835 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17814 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17808);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[4] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[3] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5894 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[3]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[9] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5377 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5377));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5926 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5485 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5485));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5345 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5345));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5890 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5926 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5892);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17821 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5894 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5890);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[6] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5905 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5909 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5916 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5909);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[7] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17945 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5452 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5452 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17945) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10862 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10862 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5924 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[15]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17828 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5916 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5924);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17811 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17821 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17828);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17829 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17811) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17835)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17829);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6374 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[28] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6262 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6262 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[29] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17952 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17952;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6364 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6364;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6474 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6474;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[31] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[31];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[31];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6249 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6249;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17959 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17959;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6462 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6462;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[34] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[34];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6235 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[33] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[33];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6235 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6349 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6349;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6158 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6158;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__44 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[0] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__44;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[44] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[44];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6412 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[43] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[43];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[42] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[42];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[41] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[41];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[40] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[40];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[39] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[39];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[38] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[38];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[37] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[37];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[36] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[36];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[35] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[35];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6436 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6256 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6366 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6256);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6476 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6436) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6366);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6412) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6476;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6198 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6294 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6439 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6223 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6439);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6334 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6294) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6223);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6198) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6334;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[46] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[46];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6186 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[45] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[45];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6393 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6213 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6324 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6213);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6434 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6393) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6324);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6186) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6434;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6303 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6253 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6395 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6178 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6395);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6292 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6253) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6178);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6303) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6292;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[47] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[47];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6402 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6210 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6244 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6357 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6244);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6466 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6357);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6251 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6210) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6466);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6402) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6251;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023 & b_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023) & a_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[48] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[48];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6288 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6354 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6384 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6168 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6384);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6280 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6168);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6391 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6354) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6280);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6288) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6391;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[49] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[49];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6166 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6200 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6199 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6200);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6314 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6199);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6423 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6314);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6207 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6166) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6423);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10745 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6207;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10745;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6311 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6344 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386) & (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6454 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6344);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6239 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6454);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6352 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6311) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6239);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6352;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6339 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6208 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6339) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6208;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6464 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6449 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6464) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6449;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6440 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6351 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6440) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6351;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6414 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6226 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6226 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6414) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6226) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6315 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6478 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6404 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6188 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6478) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6404);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6315) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6188;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17752 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17767 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17752 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17776 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17754 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17776;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17746 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17746 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17754) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17746) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17767));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6214 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6447 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6214 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6447;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6187 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6328 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6328 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6187) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6328) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6839 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6764 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6839) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6764);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7345 = (N8667 & N8664) | ((!N8667) & N8662);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225 = !(N9669 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7345);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7199 = (N8667 & N8692) | ((!N8667) & N8690);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265 = !(N9665 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7199);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6782 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6811 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6831 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6851 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6811) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6831);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6782) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17637 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 = !N8835;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7216 = (N8703 & N8728) | ((!N8703) & N8726);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298 = !(N9669 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7216);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7236 = (N8667 & N8685) | ((!N8667) & N8683);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339 = !(N9665 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7236);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6785 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6807 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6826 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6848 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6807) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6826);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6836 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6856 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6783 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6836) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6856);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6772 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6848) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6783);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6801 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6785 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6772);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6769 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6790 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6812 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6769) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6790);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6798 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6819 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6840 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6798) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6819);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6815 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6812) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6840);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6827 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6849 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6775 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6827) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6849);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6760 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10869 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6760);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6804 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10869;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6855 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6775) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6804);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6843 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6815 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6855);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[0] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6801)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6843);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 = !N9037;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7273 = (N8667 & N8671) | ((!N8667) & N8669);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246 = !(N9667 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7273);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294 = (N8696 & N8700) | ((!N8696) & N8698);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287 = !(N9665 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17644 = (N8667 & N8678) | ((!N8667) & N8785);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7319 = !(N9668 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17644);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7331 = (N8696 & N8735) | ((!N8696) & N8733);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359 = !(N9667 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7331);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7319));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6842 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6834 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6842);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6777 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6797 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6818 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6797);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6806 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6825 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6847 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6825);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6800 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6818 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6847);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[1] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6834) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6800);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243 = !N8621;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221 = N8696 & N8726;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221 & N9666);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242 = N8696 & N8785;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242 & N9669);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316 = N8696 & N8662;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316 & N9666);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335 = N8669 & N8803;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335 & N9668);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263 = N8683 & N8803;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263 & N9666);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284 = N8733 & N8981;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284 & N9668);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357 = N8690 & N8738;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351 = !(N9663 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7781 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7323 = (N8703 & N8707) | ((!N8703) & N8692);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277 = !((N9668 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7323) | ((!N9668) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7360 = (N8703 & N8714) | ((!N8703) & N8685);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313 = !((N9667 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7360) | ((!N9667) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7211 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10715 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10721 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7252 = N8773 & N8775;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202 = !((N9669 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7252) | ((!N9669) & N8467));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17664 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17618 = !(N8785 & (!N8667));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17642 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17618 & N8643) | N8641);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17974 = !N8835;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17974;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17631 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17642 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17628 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17660 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17638 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17660 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17632 = !((N8652 & N8650) | N8641);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17626 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17649 = !(N9667 | N8657);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17648 = !((N8472 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17632) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17649);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17631 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17648);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7695 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7229 = (N8703 & N8721) | ((!N8703) & N8671);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349 = !((N9668 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7229) | ((!N9668) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7267 = (N8738 & N8749) | ((!N8738) & N8678);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7219 = !((N9666 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7267) | ((!N9666) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17655 = (N8703 & N8770) | ((!N8703) & N8735);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7240 = !((N9667 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17655) | ((!N9667) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7240) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7219));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7304 = (N8738 & N8756) | ((!N8738) & N8664);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7255 = !((N9666 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7304) | ((!N9666) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7255));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7340 = (N8738 & N8742) | ((!N8738) & N8728);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7292 = !((N9669 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7340) | ((!N9669) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7292));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7209 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7209));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7798 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7742 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7781) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7695) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7798);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204 = !(N8467 & N9663);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558 = !rm[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581 = !rm[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8 = (rm[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582 = !rm[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5 = (rm[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309 & b_sign) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309) & a_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6 = (rm[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7640 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7524 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N626 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N627 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N626 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7530 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7524 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N627;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7530 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7603 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7606 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260)) | (!N8812);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54 = (N8621 & N8625) | ((!N8621) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7606);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7625 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[2])) | (!N8457);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__53 = (N8621 & N8454) | ((!N8621) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7647 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__53) | (N8267 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7625);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N639 = ((!N6997) & (!N8274)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7661 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N639 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7647;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7661;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10790 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10790;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7670 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7208 = (N8738 & N7476) | ((!N8738) & N8761);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7327 = !((N9665 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7208) | ((!N9665) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7342 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7327));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7247 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7342) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7247));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7670) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8317 = !((rm[0] & rm[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N652 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8339 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N652 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8317) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7961 = !a_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10851 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10851;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7961) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7950 = !a_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7950) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[0] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7980 = !a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7980 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7945 = !a_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7945) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7970 = !a_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8025 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8024 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8025);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8021 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[3]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8024);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7976 = !a_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7976 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7941 = !a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7941) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8015 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[1]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8021));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7737 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7721 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7737 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7768 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7721);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7797 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7768);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7667 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7797 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7667);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17979 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[23] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17979;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N642 = !((N7476 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[23]) | N7472);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62 = !(N7364 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N642);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70 = N6992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4317 = ((a_exp[0] & a_exp[1]) & a_exp[7]) & a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4321 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4317 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4321);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4354 = !(a_man[8] | a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4352 = ((a_man[6] | a_man[4]) | a_man[5]) | a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4357 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4354) | a_man[10]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4352) | a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4377 = !(a_man[22] | a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4369 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4379 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4373 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4369 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4379);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4340 = !(a_man[20] | a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10761 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4377 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4373) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4340);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4346 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338) | a_man[0]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10761) | a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4357 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4346);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4412 = ((b_exp[0] & b_exp[1]) & b_exp[7]) & b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4416 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4412 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4416);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4447 = ((b_man[6] | b_man[4]) | b_man[5]) | b_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4437 = ((b_man[10] | b_man[8]) | b_man[9]) | b_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4454 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4462 = !(b_man[0] | b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4464 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4474 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4468 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4464 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4474);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10769 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4462) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4447 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4437) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4454) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10769;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10775 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4525 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10775);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4525;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8363 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70 | N9673;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933, fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8075} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206} + {1'B0, N7705};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[23] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8075;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8075 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243) ^ N7719;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8086 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8086;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8070 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8112 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8070;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8094 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109, fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088} = {1'B0, N9665} + {1'B0, N7727};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110 = !(N7682 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071, fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517} = {1'B0, N8803} + {1'B0, N7735};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541, fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272} + {1'B0, N7713};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529 = N7719 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8038 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090 = !(N7682 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8066 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8106 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8066);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8038) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8106);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17480 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048 & N7208) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048) & N7210));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17485 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17480);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8059 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8059) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8067 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8084 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8084) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8067);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17458 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8100 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8118 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8118) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8100);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8057 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8037 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048 & N7327) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048) & N7325);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17466 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8111 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[6] = N7317 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8082 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8082;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17475 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17470 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17458 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17466) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17475);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17493 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[5] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17483 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17493 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8058 = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17489 = ((!N7358) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048)) | ((!N7354) & (!N7356));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17456 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17489);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17463 = !(N7090 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17456);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17470 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17485) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17463);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71;
assign x[22] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8363) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7775 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7717 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7672 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7775) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7717) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7804 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7804;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10843 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7672 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10843;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7025 = !(b_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8461 = !((N9673 & N6809) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8461) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[21]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7710 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7795 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7758 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7710) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7795) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7713 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7713;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10836 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7758 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10836;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6966 = !(b_man[20] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8435 = !((N9673 & N6802) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8435) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[20]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7694 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7679 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7694 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7679;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7042 = !(b_man[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8407 = (N9671 & N6729) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[19] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8407) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7668 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7773 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7668) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7695) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7731 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7773 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7731;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6984 = !(b_man[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6984 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8379 = (N9671 & N6722) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[18] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8379) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7755 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10829 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7755) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7775) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10829;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7060 = !(b_man[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7060 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8353 = !((N9673 & N6795) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8353) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[17]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7691 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7791 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7691) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7710) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7684 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7791 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7684;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7000 = !(b_man[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7000 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8451 = (N9671 & N6715) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[16] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8451) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7806 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7806;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7076 = !(b_man[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8424 = (N9671 & N6708) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[15] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8424) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7716 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7781 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7716;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7016 = !(b_man[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8394 = (N9671 & N6701) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[14] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8394) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10822 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7717 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7804);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[13] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10822;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7092 = !(b_man[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8368 = !((N9673 & N6788) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8368) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[13]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10815 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7795 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7713);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[12] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10815;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7035 = !(b_man[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7035 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8466 = !((N9673 & N6781) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8466) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[12]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10808 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10808;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6977 = !(b_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8440 = !((N9673 & N6774) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8440) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[11]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10801 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7668 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[10] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10801;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7054 = !(b_man[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7054 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8412 = !((N9673 & N6767) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8412) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7675 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7755 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7675;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6995 = !(b_man[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6995 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8384 = (N9671 & N6694) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[9] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8384) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10794 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7691 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10794;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7071 = !(b_man[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8358 = !((N9673 & N6760) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8358) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7667) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7011 = !(b_man[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7011 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8456 = (N9671 & N6687) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8456) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7086 = !(b_man[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7086 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8429 = !((N9673 & N6753) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8429) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7028 = !(b_man[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7028 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8400 = (N9671 & N6680) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8400) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6969 = !(b_man[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6969 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8373 = (N9671 & N6673) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8373) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7045 = !(b_man[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7045 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8346 = !((N9673 & N6746) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8346) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[3]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6987 = !(b_man[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6987 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8445 = !((N9673 & N6739) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8445) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7064 = !(b_man[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7064) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8417 = (N9671 & N6666) | ((!N9671) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70);
assign x[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8417) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7004 = !(b_man[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[0] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7004 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8388 = !((N9673 & N6732) | ((!N9673) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70));
assign x[0] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8388) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8253 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296 = !(N6821 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71;
assign x[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[7]));
assign x[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[6]));
assign x[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[5]));
assign x[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[4]));
assign x[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[3]));
assign x[25] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8276 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[1];
assign x[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8276));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8243 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4) | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N651 = !(((!N6999) & (!N6997)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[0] = N6821 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N651;
assign x[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17966 = a_sign | b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N645 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6) | (a_sign & b_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6958 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__66 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N645 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6958);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7050 = !(b_sign | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7017 = !a_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N710 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7050) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7182 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N710) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63) & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__66));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7185 = !((N6959 & N6955) | ((!N6959) & N6957));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7191 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63 | fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706);
assign x[31] = !((N6624 & fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7185) | ((!N6624) & N6622));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[30] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[34] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[35] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[36] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[38] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[39] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[40] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[41] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  v7XxSQ3arBw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



