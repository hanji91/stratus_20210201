/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:25:18 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895;
wire N5143,N5150,N5157,N5164,N5171,N5178,N5185 
	,N5192,N5199,N5206,N5213,N5220,N5227,N5234,N5241 
	,N5248,N5255,N5262,N5269,N5276,N5283,N5295,N5354 
	,N5356,N5592,N5605,N5607,N5631,N5633,N5712,N5717 
	,N5967,N5998,N6004,N6029,N6042,N6048,N6069,N6071 
	,N6079,N6091,N6093,N6099,N6101,N6111,N6119,N6137 
	,N6171,N6182,N6563,N6570,N6572,N6873,N6875,N6880 
	,N6882,N6887,N6889,N6894,N6896,N6899,N6901,N6903 
	,N6908,N6925,N7051,N7053,N7058,N7060,N7063,N7209 
	,N7216,N7318,N7325,N7348,N7368,N7375,N7382,N7389 
	,N7396,N7440,N7536,N7540,N7577,N7604,N7608,N7714 
	,N7720,N7722,N7724,N7727,N7729,N7731,N7998,N8000 
	,N8191,N8192,N8193,N8194;
reg x_reg_15__retimed_I4479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4479_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996;
	end
assign N8000 = x_reg_15__retimed_I4479_QOUT;
reg x_reg_15__retimed_I4478_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4478_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000;
	end
assign N7998 = x_reg_15__retimed_I4478_QOUT;
reg x_reg_15__retimed_I4366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4366_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046;
	end
assign N7731 = x_reg_15__retimed_I4366_QOUT;
reg x_reg_15__retimed_I4365_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4365_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061;
	end
assign N7729 = x_reg_15__retimed_I4365_QOUT;
reg x_reg_15__retimed_I4364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4364_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086;
	end
assign N7727 = x_reg_15__retimed_I4364_QOUT;
reg x_reg_15__retimed_I4363_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4363_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997;
	end
assign N7724 = x_reg_15__retimed_I4363_QOUT;
reg x_reg_15__retimed_I4362_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4362_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070;
	end
assign N7722 = x_reg_15__retimed_I4362_QOUT;
reg x_reg_15__retimed_I4361_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4361_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011;
	end
assign N7720 = x_reg_15__retimed_I4361_QOUT;
reg x_reg_15__retimed_I4360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4360_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032;
	end
assign N7714 = x_reg_15__retimed_I4360_QOUT;
reg x_reg_15__retimed_I4344_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4344_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049;
	end
assign N7608 = x_reg_15__retimed_I4344_QOUT;
reg x_reg_15__retimed_I4342_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4342_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078;
	end
assign N7604 = x_reg_15__retimed_I4342_QOUT;
reg x_reg_15__retimed_I4334_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4334_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065;
	end
assign N7577 = x_reg_15__retimed_I4334_QOUT;
reg x_reg_15__retimed_I4331_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4331_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082;
	end
assign N7540 = x_reg_15__retimed_I4331_QOUT;
reg x_reg_15__retimed_I4329_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4329_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014;
	end
assign N7536 = x_reg_15__retimed_I4329_QOUT;
reg x_reg_15__retimed_I4313_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4313_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655;
	end
assign N7440 = x_reg_15__retimed_I4313_QOUT;
reg x_reg_15__retimed_I4297_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4297_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3];
	end
assign N7396 = x_reg_15__retimed_I4297_QOUT;
reg x_reg_15__retimed_I4294_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4294_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4];
	end
assign N7389 = x_reg_15__retimed_I4294_QOUT;
reg x_reg_15__retimed_I4291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4291_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N7382 = x_reg_15__retimed_I4291_QOUT;
reg x_reg_15__retimed_I4288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4288_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N7375 = x_reg_15__retimed_I4288_QOUT;
reg x_reg_15__retimed_I4285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4285_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N7368 = x_reg_15__retimed_I4285_QOUT;
reg x_reg_15__retimed_I4277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4277_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
	end
assign N7348 = x_reg_15__retimed_I4277_QOUT;
reg x_reg_15__retimed_I4273_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4273_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
	end
assign N7325 = x_reg_15__retimed_I4273_QOUT;
reg x_reg_15__retimed_I4270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4270_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6];
	end
assign N7318 = x_reg_15__retimed_I4270_QOUT;
reg x_reg_15__retimed_I4238_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4238_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8];
	end
assign N7216 = x_reg_15__retimed_I4238_QOUT;
reg x_reg_15__retimed_I4235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4235_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7];
	end
assign N7209 = x_reg_15__retimed_I4235_QOUT;
reg x_reg_15__retimed_I4188_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4188_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4;
	end
assign N7063 = x_reg_15__retimed_I4188_QOUT;
reg x_reg_15__retimed_I4187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4187_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17];
	end
assign N7060 = x_reg_15__retimed_I4187_QOUT;
reg x_reg_15__retimed_I4186_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4186_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
	end
assign N7058 = x_reg_15__retimed_I4186_QOUT;
reg x_reg_15__retimed_I4184_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4184_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18];
	end
assign N7053 = x_reg_15__retimed_I4184_QOUT;
reg x_reg_15__retimed_I4183_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4183_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10];
	end
assign N7051 = x_reg_15__retimed_I4183_QOUT;
reg x_reg_15__retimed_I4139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4139_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638;
	end
assign N6925 = x_reg_15__retimed_I4139_QOUT;
reg x_reg_15__retimed_I4132_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4132_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43;
	end
assign N6908 = x_reg_15__retimed_I4132_QOUT;
reg x_reg_15__retimed_I4130_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4130_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
	end
assign N6903 = x_reg_15__retimed_I4130_QOUT;
reg x_reg_15__retimed_I4129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4129_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635;
	end
assign N6901 = x_reg_15__retimed_I4129_QOUT;
reg x_reg_15__retimed_I4128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4128_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N6899 = x_reg_15__retimed_I4128_QOUT;
reg x_reg_15__retimed_I4127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4127_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21];
	end
assign N6896 = x_reg_15__retimed_I4127_QOUT;
reg x_reg_15__retimed_I4126_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4126_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
	end
assign N6894 = x_reg_15__retimed_I4126_QOUT;
reg x_reg_15__retimed_I4124_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4124_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22];
	end
assign N6889 = x_reg_15__retimed_I4124_QOUT;
reg x_reg_15__retimed_I4123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4123_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14];
	end
assign N6887 = x_reg_15__retimed_I4123_QOUT;
reg x_reg_15__retimed_I4121_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4121_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20];
	end
assign N6882 = x_reg_15__retimed_I4121_QOUT;
reg x_reg_15__retimed_I4120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4120_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12];
	end
assign N6880 = x_reg_15__retimed_I4120_QOUT;
reg x_reg_15__retimed_I4118_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4118_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19];
	end
assign N6875 = x_reg_15__retimed_I4118_QOUT;
reg x_reg_15__retimed_I4117_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4117_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11];
	end
assign N6873 = x_reg_15__retimed_I4117_QOUT;
reg x_reg_15__retimed_I4000_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4000_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23];
	end
assign N6572 = x_reg_15__retimed_I4000_QOUT;
reg x_reg_15__retimed_I3999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3999_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15];
	end
assign N6570 = x_reg_15__retimed_I3999_QOUT;
reg x_reg_15__retimed_I3996_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3996_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16];
	end
assign N6563 = x_reg_15__retimed_I3996_QOUT;
reg x_reg_15__retimed_I3848_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3848_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0];
	end
assign N6182 = x_reg_15__retimed_I3848_QOUT;
reg x_reg_15__retimed_I3844_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3844_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
	end
assign N6171 = x_reg_15__retimed_I3844_QOUT;
reg x_reg_15__retimed_I3832_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3832_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918;
	end
assign N6137 = x_reg_15__retimed_I3832_QOUT;
reg x_reg_15__retimed_I3825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3825_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944;
	end
assign N6119 = x_reg_15__retimed_I3825_QOUT;
reg x_reg_15__retimed_I3822_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3822_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911;
	end
assign N6111 = x_reg_15__retimed_I3822_QOUT;
reg x_reg_15__retimed_I3818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3818_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923;
	end
assign N6101 = x_reg_15__retimed_I3818_QOUT;
reg x_reg_15__retimed_I3817_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3817_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936;
	end
assign N6099 = x_reg_15__retimed_I3817_QOUT;
reg x_reg_15__retimed_I3815_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3815_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928;
	end
assign N6093 = x_reg_15__retimed_I3815_QOUT;
reg x_reg_15__retimed_I3814_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3814_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
	end
assign N6091 = x_reg_15__retimed_I3814_QOUT;
reg x_reg_15__retimed_I3809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3809_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
	end
assign N6079 = x_reg_15__retimed_I3809_QOUT;
reg x_reg_15__retimed_I3806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3806_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24];
	end
assign N6071 = x_reg_15__retimed_I3806_QOUT;
reg x_reg_15__retimed_I3805_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3805_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
	end
assign N6069 = x_reg_15__retimed_I3805_QOUT;
reg x_reg_15__retimed_I3798_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3798_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901;
	end
assign N6048 = x_reg_15__retimed_I3798_QOUT;
reg x_reg_15__retimed_I3796_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3796_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921;
	end
assign N6042 = x_reg_15__retimed_I3796_QOUT;
reg x_reg_15__retimed_I3791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3791_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883;
	end
assign N6029 = x_reg_15__retimed_I3791_QOUT;
reg x_reg_15__retimed_I3783_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3783_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908;
	end
assign N6004 = x_reg_15__retimed_I3783_QOUT;
reg x_reg_15__retimed_I3781_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3781_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929;
	end
assign N5998 = x_reg_15__retimed_I3781_QOUT;
reg x_reg_15__retimed_I3768_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3768_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018;
	end
assign N5967 = x_reg_15__retimed_I3768_QOUT;
reg x_reg_23__retimed_I3675_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3675_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650;
	end
assign N5717 = x_reg_23__retimed_I3675_QOUT;
reg x_reg_22__retimed_I3673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3673_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111;
	end
assign N5712 = x_reg_22__retimed_I3673_QOUT;
reg x_reg_31__retimed_I3668_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3668_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6;
	end
assign N5633 = x_reg_31__retimed_I3668_QOUT;
reg x_reg_31__retimed_I3667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3667_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
	end
assign N5631 = x_reg_31__retimed_I3667_QOUT;
reg x_reg_23__retimed_I3659_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3659_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17;
	end
assign N5607 = x_reg_23__retimed_I3659_QOUT;
reg x_reg_23__retimed_I3658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3658_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12;
	end
assign N5605 = x_reg_23__retimed_I3658_QOUT;
reg x_reg_15__retimed_I3656_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3656_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
	end
assign N5592 = x_reg_15__retimed_I3656_QOUT;
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4575 (.Y(N8191), .A(N5592));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4576 (.Y(N8192), .A(N8191));
reg x_reg_31__retimed_I3561_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3561_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282;
	end
assign N5356 = x_reg_31__retimed_I3561_QOUT;
reg x_reg_31__retimed_I3560_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3560_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291;
	end
assign N5354 = x_reg_31__retimed_I3560_QOUT;
reg x_reg_15__retimed_I3535_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3535_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15];
	end
assign N5295 = x_reg_15__retimed_I3535_QOUT;
reg x_reg_0__retimed_I3530_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3530_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0];
	end
assign N5283 = x_reg_0__retimed_I3530_QOUT;
reg x_reg_1__retimed_I3527_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I3527_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1];
	end
assign N5276 = x_reg_1__retimed_I3527_QOUT;
reg x_reg_2__retimed_I3524_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I3524_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2];
	end
assign N5269 = x_reg_2__retimed_I3524_QOUT;
reg x_reg_3__retimed_I3521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I3521_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3];
	end
assign N5262 = x_reg_3__retimed_I3521_QOUT;
reg x_reg_4__retimed_I3518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I3518_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4];
	end
assign N5255 = x_reg_4__retimed_I3518_QOUT;
reg x_reg_5__retimed_I3515_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I3515_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5];
	end
assign N5248 = x_reg_5__retimed_I3515_QOUT;
reg x_reg_6__retimed_I3512_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3512_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6];
	end
assign N5241 = x_reg_6__retimed_I3512_QOUT;
reg x_reg_7__retimed_I3509_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3509_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7];
	end
assign N5234 = x_reg_7__retimed_I3509_QOUT;
reg x_reg_8__retimed_I3506_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3506_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8];
	end
assign N5227 = x_reg_8__retimed_I3506_QOUT;
reg x_reg_9__retimed_I3503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3503_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9];
	end
assign N5220 = x_reg_9__retimed_I3503_QOUT;
reg x_reg_10__retimed_I3500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3500_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10];
	end
assign N5213 = x_reg_10__retimed_I3500_QOUT;
reg x_reg_11__retimed_I3497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3497_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11];
	end
assign N5206 = x_reg_11__retimed_I3497_QOUT;
reg x_reg_12__retimed_I3494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3494_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12];
	end
assign N5199 = x_reg_12__retimed_I3494_QOUT;
reg x_reg_13__retimed_I3491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3491_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13];
	end
assign N5192 = x_reg_13__retimed_I3491_QOUT;
reg x_reg_14__retimed_I3488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3488_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14];
	end
assign N5185 = x_reg_14__retimed_I3488_QOUT;
reg x_reg_16__retimed_I3485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3485_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16];
	end
assign N5178 = x_reg_16__retimed_I3485_QOUT;
reg x_reg_17__retimed_I3482_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3482_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17];
	end
assign N5171 = x_reg_17__retimed_I3482_QOUT;
reg x_reg_18__retimed_I3479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3479_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18];
	end
assign N5164 = x_reg_18__retimed_I3479_QOUT;
reg x_reg_19__retimed_I3476_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I3476_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19];
	end
assign N5157 = x_reg_19__retimed_I3476_QOUT;
reg x_reg_20__retimed_I3473_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I3473_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20];
	end
assign N5150 = x_reg_20__retimed_I3473_QOUT;
reg x_reg_21__retimed_I3470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I3470_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21];
	end
assign N5143 = x_reg_21__retimed_I3470_QOUT;
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I0 (.Y(bdw_enable), .A(astall));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132), .A(a_exp[0]), .B(a_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I2 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I3 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834), .A(a_exp[7]), .B(a_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I6 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I7 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155), .A(a_man[10]), .B(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I8 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174), .A(a_man[6]), .B(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I9 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163), .A(a_man[8]), .B(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I10 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183), .A(a_man[4]), .B(a_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I11 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I12 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I13 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I14 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I15 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I16 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[7]), .D(b_exp[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I17 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559), .A(b_exp[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I18 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I19 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I20 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I21 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I22 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I23 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232), .A(b_man[10]), .B(b_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I24 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251), .A(b_man[6]), .B(b_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I25 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240), .A(b_man[8]), .B(b_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I26 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260), .A(b_man[4]), .B(b_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I27 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I28 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I29 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I30 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I31 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I32 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I33 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I34 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I35 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
OR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I36 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I37 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563), .A(b_exp[7]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I38 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408), .A(a_exp[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I39 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562), .A(b_exp[6]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I40 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376), .A(a_exp[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I41 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561), .A(b_exp[5]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I42 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418), .A(a_exp[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I43 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560), .A(b_exp[4]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I44 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386), .A(a_exp[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I45 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360), .A(a_exp[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I46 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558), .A(b_exp[2]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I47 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396), .A(a_exp[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I48 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733), .A(a_exp[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I49 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557), .A(b_exp[1]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I50 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730), .A(a_exp[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I51 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I52 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556), .A(b_exp[0]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I53 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I54 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372), .A(a_exp[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I55 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I56 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380), .A(a_exp[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I57 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I58 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I59 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377), .A(a_exp[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I60 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I61 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417), .A(a_exp[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I62 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I63 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382), .A(a_exp[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I64 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I65 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357), .A(a_exp[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I66 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I67 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393), .A(a_exp[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I68 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I69 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I70 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I71 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556), .B(a_exp[0]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I72 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I73 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I74 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I75 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I76 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I77 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I78 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I79 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I80 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I81 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520), .A(a_man[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I82 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538), .A(b_man[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I83 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607), .A(a_man[21]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I84 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I85 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541), .A(a_man[20]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I86 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I87 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I88 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I89 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473), .A(a_man[19]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I90 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I91 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561), .A(a_man[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I92 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I93 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I94 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494), .A(a_man[17]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I95 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I96 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578), .A(a_man[16]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I97 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I98 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I99 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552), .A(a_man[11]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I101 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484), .A(a_man[10]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I104 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I105 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570), .A(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I106 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I107 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516), .A(a_man[15]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I108 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I109 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598), .A(a_man[14]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I110 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531), .A(a_man[13]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I114 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468), .A(a_man[12]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507), .A(a_man[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588), .A(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I123 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524), .A(a_man[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I124 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I125 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I126 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610), .A(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I127 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I128 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543), .A(a_man[4]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I129 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I130 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I131 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I132 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478), .A(a_man[3]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I133 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I134 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564), .A(a_man[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I135 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I136 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I137 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504), .A(b_man[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I138 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497), .A(a_man[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I139 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I140 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497));
OAI31X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I141 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504), .A1(a_man[0]), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I142 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I143 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I144 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I145 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I146 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I147 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I148 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I149 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I150 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I151 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I152 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I153 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I154 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I155 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I156 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I157 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I158 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I159 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I160 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I161 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I162 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I163 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I164 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I165 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I166 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I167 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I168 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I169 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I170 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I171 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I172 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I173 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I174 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I175 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I176 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I177 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I178 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I179 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I180 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536), .B0(b_man[22]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I181 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I182 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I183 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I184 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575));
CLKINVX6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I185 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I186 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .A(a_man[15]), .B(b_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I187 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I188 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I189 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I190 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340), .A(b_exp[7]), .B(b_exp[5]), .C(b_exp[6]), .D(b_exp[4]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I191 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I192 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I193 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16));
BUFX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I194 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I195 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I196 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I197 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I198 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I199 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I200 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I201 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I202 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I203 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I204 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I205 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I206 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I207 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I208 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I209 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I210 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
OAI211X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I211 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I212 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I213 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I214 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I215 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I216 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I217 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I218 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I219 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I220 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I221 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I222 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I223 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I224 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I225 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .A(b_man[20]), .B(a_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I226 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .A(b_man[19]), .B(a_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I227 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0]), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I228 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I229 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I230 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I231 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I232 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I233 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I234 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I235 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I236 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I237 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I238 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I239 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I240 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I241 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I242 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I243 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I244 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I245 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I246 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I247 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I248 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I249 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I250 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I251 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I252 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I253 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I254 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I255 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I256 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .A(a_man[14]), .B(b_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I257 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I258 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .A(b_man[14]), .B(a_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I259 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I260 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I261 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I262 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I263 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I264 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I265 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I266 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I267 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I269 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I270 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I271 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I272 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I273 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I274 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .A(a_man[13]), .B(b_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I275 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .A(b_man[13]), .B(a_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I276 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I277 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I278 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I279 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I280 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I281 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I282 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I283 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I284 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I285 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I286 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I287 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I288 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .A(a_man[12]), .B(b_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I289 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I290 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I291 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I292 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I293 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I294 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I295 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I296 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I297 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I298 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I299 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I300 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I301 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .A(a_man[11]), .B(b_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I302 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .A(b_man[11]), .B(a_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I303 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I304 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I305 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I306 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I307 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I308 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I309 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I310 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I311 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I312 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I313 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I314 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I315 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I316 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .A(a_man[10]), .B(b_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I317 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I318 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I319 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I320 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I321 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I322 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I323 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I324 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I325 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I326 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I327 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I328 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I329 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .A(a_man[9]), .B(b_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I330 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I331 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I332 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I333 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I334 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I335 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I336 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I337 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I338 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I339 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I340 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I341 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I342 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .A(a_man[8]), .B(b_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I343 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I344 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I345 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I346 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I347 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I348 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I349 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I350 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I351 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I352 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I353 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I354 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .A(a_man[7]), .B(b_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I355 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I356 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I357 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I358 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I359 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I360 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I361 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I362 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I363 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I364 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I365 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I366 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I367 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I368 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .A(a_man[6]), .B(b_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I369 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I370 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I371 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I372 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I373 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I374 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I375 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I376 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I377 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I378 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660), .A(a_man[5]), .B(b_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I379 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I380 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I381 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I382 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I383 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I384 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I385 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I386 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I387 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I388 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659), .A(a_man[4]), .B(b_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I390 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .A(b_man[4]), .B(a_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I391 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I392 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I393 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I394 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I396 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I397 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I398 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I399 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .A(a_man[3]), .B(b_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I400 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .A(b_man[3]), .B(a_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I401 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I402 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I403 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I404 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I407 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I409 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I412 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I413 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I415 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I416 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I417 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I418 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I419 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I420 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I421 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656), .A(a_man[1]), .B(b_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I422 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I423 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I424 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I425 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I427 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I428 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I429 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I430 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I431 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I432 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .A(a_man[0]), .B(b_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I433 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .A(b_man[0]), .B(a_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I434 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I435 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I436 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I437 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I438 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I439 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I440 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I441 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I442 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I443 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I444 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I445 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I446 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I447 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I448 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I449 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I450 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I451 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I452 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I453 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I454 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I455 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I456 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I457 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I458 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I459 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I460 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I461 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I462 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I463 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I464 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I465 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I466 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I467 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I468 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I469 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I470 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I471 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I472 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I473 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I474 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I475 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I476 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I477 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I478 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I479 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I480 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I481 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I482 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I483 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I484 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I485 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I486 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I487 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I488 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I489 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I490 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I491 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I492 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I493 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I494 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I495 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I496 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I497 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I498 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I499 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I500 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I501 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I502 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I503 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I504 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I505 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I506 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I507 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I508 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I509 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I510 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I511 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I512 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I513 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I514 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I515 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I516 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I517 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I518 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I519 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I520 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I521 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I522 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I523 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I524 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I525 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436));
NAND2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I526 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I527 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I528 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I529 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I530 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I531 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I532 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I533 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I534 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I535 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I536 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I537 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I538 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I539 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I540 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I541 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I542 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I543 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I544 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I545 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I546 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I547 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I548 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I549 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I550 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I551 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I552 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I553 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I554 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I555 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I556 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I557 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I558 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I559 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I560 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I561 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I562 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I563 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I564 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .A(a_man[16]), .B(b_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I565 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I566 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I567 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I568 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I569 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I570 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I571 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I572 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I573 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I574 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I575 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I576 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I577 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I578 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I579 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I580 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I581 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I582 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I583 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I584 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I585 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I586 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I587 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I588 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I589 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I590 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I591 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I592 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I593 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I594 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I595 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I596 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I597 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I598 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I599 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I600 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I601 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .A(a_man[22]), .B(b_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I602 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I603 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I604 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I605 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .A(a_man[21]), .B(b_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I606 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I607 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I608 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I609 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I610 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .A(a_man[20]), .B(b_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I611 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I612 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I613 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I614 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .A(a_man[19]), .B(b_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I615 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I616 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I617 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I618 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I619 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .A(a_man[18]), .B(b_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I620 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I621 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I622 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I623 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .A(a_man[17]), .B(b_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I624 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I625 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I626 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I627 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I628 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I629 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I630 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I631 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I632 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I633 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I634 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I635 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I636 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I637 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I638 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I639 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I640 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I641 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I642 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I643 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823));
OAI31X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I644 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I645 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I646 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I647 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I648 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I649 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I650 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I651 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I652 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I653 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I654 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I655 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I656 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I657 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I658 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I659 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I660 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I661 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I662 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I663 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I664 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I665 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I666 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I667 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010), .A(N7720), .B(N7729));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I668 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I669 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I670 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I671 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I672 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I673 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I674 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I675 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I676 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I677 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I678 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I679 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I680 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I681 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I682 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I683 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I684 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I685 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I686 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I687 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I688 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I689 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I690 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I691 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I692 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I693 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I694 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I695 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I696 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I697 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I698 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I699 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I700 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031), .A0(N7729), .A1(N7608), .B0(N7604));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I701 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010), .A1(N7577), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I702 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919), .A(N6171), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I703 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I704 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I705 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I706 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I707 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I708 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I709 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I710 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I711 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I712 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I713 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I714 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I715 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I716 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I717 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I718 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I719 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I720 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I721 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I722 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I723 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I724 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I725 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I726 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I727 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I728 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I729 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I730 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I731 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074), .A0(N7729), .A1(N7731), .B0(N7727));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I732 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010), .A1(N7714), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I733 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I734 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I735 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I736 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I737 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I738 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I739 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360), .A0(N7536), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010), .B0(N7540));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I740 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I741 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4577 (.Y(N8193), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4578 (.Y(N8194), .A(N8193));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I742 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I743 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039), .A(N7998), .B(N8000));
NAND2BX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I744 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I745 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I746 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I747 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061));
AO21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I748 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439), .A0(N7722), .A1(N7720), .B0(N7724));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I749 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I750 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I751 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809), .B(N7389));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I752 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I753 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328), .A(N6880), .B(N6882), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I754 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I755 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809), .B(N7396));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I756 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457), .A(N6873), .B(N6875), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I757 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I758 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I759 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I760 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I761 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I762 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I763 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392), .A(N7368), .B(N7216), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I764 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307), .A(N6563), .B(N6071), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I765 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I766 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808), .B(N7209));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I767 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436), .A(N6570), .B(N6572), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I768 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I769 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I770 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I771 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809), .B(N7375));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I772 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420), .A(N7051), .B(N7053), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I773 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I774 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383), .A(N7382), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I775 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386), .A(N7058), .B(N7060), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I776 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I777 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I778 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808), .B(N7318));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I779 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400), .A(N6887), .B(N6889), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I780 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I781 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808), .B(N7325));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I782 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365), .A(N6894), .B(N6896), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I783 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I784 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I785 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I786 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I787 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I788 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I789 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I790 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439), .B(N7368));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I791 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349), .A(N7216), .B(N6563), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I792 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I793 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I794 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I795 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I796 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I797 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I798 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441), .A(N7318), .B(N6887), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I799 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I800 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405), .A(N7325), .B(N6894), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I801 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I802 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I803 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I804 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I805 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371), .A(N7389), .B(N6880), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I806 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I807 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334), .A(N7396), .B(N6873), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I808 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I809 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I810 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315), .A(N7209), .B(N6570), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I811 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I812 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I813 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I814 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I815 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I816 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I817 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297), .A(N7375), .B(N7051), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I818 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I819 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I820 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I821 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I822 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I823 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I824 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I825 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I826 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I827 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I828 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427), .A(N7382), .B(N7058), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I829 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I830 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I831 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I832 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I833 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I834 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I835 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I836 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I837 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I838 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I839 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I840 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I841 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I842 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I843 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I844 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I845 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I846 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I847 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I848 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I849 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I850 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I851 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I852 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I853 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I854 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I855 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I856 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I857 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I858 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I859 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I860 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I861 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I862 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I863 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I864 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I865 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734));
NAND4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I866 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I867 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I868 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I869 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I870 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I871 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I872 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I873 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I874 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I875 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362), .A0(N8194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I876 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I877 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I878 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I879 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I880 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I881 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I882 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I883 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I884 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I885 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I886 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I887 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I888 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]), .B(N6908), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I889 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I890 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I891 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48), .A(b_sign), .B(a_sign), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I892 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I893 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I894 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I895 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I896 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I897 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I898 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I899 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I900 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I901 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308), .B0(N7440));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I902 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631), .B(N7348), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I903 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I904 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633), .A(N7063), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I905 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636), .A(N6903), .B(N6901), .C(N6899), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I906 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I907 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639), .A(N6925), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54));
AOI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I908 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639));
OR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I909 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I910 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I911 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I912 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I913 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769));
NAND4BX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I914 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I915 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759));
NAND4BX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I916 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I917 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I918 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I919 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I920 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I921 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777));
XOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I922 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951), .A(N6182), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I923 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941), .A(N6182), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I924 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I925 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909), .A(N6171), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I926 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I927 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I928 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I929 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946), .A(N6137), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I930 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I931 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]), .A(a_exp[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I932 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I933 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913), .A(N6119), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439));
AOI2BB2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I934 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917), .A0N(N6137), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946));
OAI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I935 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917), .B0(N6119), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I936 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I937 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I938 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938), .A(N6111), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I939 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938));
AOI2BB2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I940 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932), .A0N(N6111), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I941 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I942 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I943 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I944 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932), .B(N6004));
OAI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I945 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905), .A0(N6004), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932), .B0(N6099), .B1(N6101));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I946 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]), .A(a_exp[6]), .B(b_exp[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I947 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I948 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I949 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905), .B(N5998));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I950 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]));
AOI2BB2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I951 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930), .A0N(N6091), .A1N(N6093), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905), .B1(N5998));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I952 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]), .A(a_exp[7]), .B(b_exp[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I953 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I954 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I955 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930), .B(N6048));
OAI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I956 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950), .A0(N6048), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930), .B0(N6079), .B1(N6042));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I957 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8]), .A(N6042), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I958 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I959 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I960 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I961 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I962 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I963 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I964 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I965 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I966 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I967 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I968 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I969 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I970 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I971 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642), .A0(N6071), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]), .B0(N6069));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I972 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .A(N6029), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I973 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9]), .A(N6042), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I974 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020), .A(N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9]));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I975 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020));
NOR2BX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I976 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .AN(N8192), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I977 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092), .A(rm[0]), .B(rm[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I978 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7), .A(rm[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I979 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I980 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I981 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I982 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A(N5712), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I983 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I984 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I985 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .A(N8192), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I986 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I987 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I988 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I989 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I990 (.Y(x[22]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I991 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I992 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[21]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[21]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I993 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I994 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I995 (.Y(x[21]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5143), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I996 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[20]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[20]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I997 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I998 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I999 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1000 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1001 (.Y(x[20]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1002 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[19]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[19]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1003 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1004 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1005 (.Y(x[19]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5157), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1006 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[18]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[18]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1007 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1008 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1009 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1010 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1011 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1012 (.Y(x[18]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5164), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1013 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[17]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[17]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1014 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1015 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1016 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1017 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1018 (.Y(x[17]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5171), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1019 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[16]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1020 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1021 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1022 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1023 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1024 (.Y(x[16]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5178), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1025 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[15]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[15]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1026 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1027 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1028 (.Y(x[15]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5295), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1029 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[14]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[14]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1030 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1031 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1032 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1033 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1034 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1035 (.Y(x[14]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5185), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1036 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[13]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[13]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1037 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1038 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1039 (.Y(x[13]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5192), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1040 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[12]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1041 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1042 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1043 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1044 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1045 (.Y(x[12]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5199), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1046 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[11]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[11]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1047 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1048 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1049 (.Y(x[11]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5206), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1050 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[10]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[10]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1051 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1052 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1053 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1054 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1055 (.Y(x[10]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5213), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1056 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[9]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[9]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1057 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1058 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1059 (.Y(x[9]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5220), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1060 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1061 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1062 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1063 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1064 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1065 (.Y(x[8]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5227), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1066 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[7]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[7]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1067 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1068 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1069 (.Y(x[7]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5234), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1070 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[6]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[6]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1071 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1072 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1073 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1074 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1075 (.Y(x[6]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5241), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1076 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[5]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[5]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1077 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1078 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1079 (.Y(x[5]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5248), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1080 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[4]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1081 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1082 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1083 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1084 (.Y(x[4]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5255), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1085 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[3]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[3]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1086 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1087 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1088 (.Y(x[3]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5262), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1089 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[2]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[2]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1090 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1091 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1092 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1093 (.Y(x[2]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5269), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1094 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[1]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1095 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1096 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1097 (.Y(x[1]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5276), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1098 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[0]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_man[0]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1099 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1101 (.Y(x[0]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141), .A1N(N5283), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .A(N5605), .B(N5607), .C(N5592), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1104 (.Y(x[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1105 (.Y(x[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1106 (.Y(x[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1107 (.Y(x[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1108 (.Y(x[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1109 (.Y(x[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1110 (.Y(x[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651), .A(N5717), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]), .A(N5605), .B(N5607), .C(N8192), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1114 (.Y(x[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895), .A(a_sign), .B(b_sign));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233), .A0(a_sign), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212), .B1(b_sign));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285), .A(N5631), .B(N5633), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1123 (.Y(x[31]), .A(N5356), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285), .S0(N5354));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[28] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  v7P4Sg/WqB0= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



